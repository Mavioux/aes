module MixColumns (
    input wire [0:127] state,
    output reg [0:127] new_state
);
    

endmodule