module MixColumn1RowInverse (
    input wire [0:31] row,
    output wire [0:7] output_row
);
    reg [0:7] a, b, c, d;

    // Multiplication with 14
    always @(row[0:7]) begin
        case (row[0:7])
            8'h0 : a[0:7] = 8'h0;
            8'h1 : a[0:7] = 8'he;
            8'h2 : a[0:7] = 8'h1c;
            8'h3 : a[0:7] = 8'h12;
            8'h4 : a[0:7] = 8'h38;
            8'h5 : a[0:7] = 8'h36;
            8'h6 : a[0:7] = 8'h24;
            8'h7 : a[0:7] = 8'h2a;
            8'h8 : a[0:7] = 8'h70;
            8'h9 : a[0:7] = 8'h7e;
            8'ha : a[0:7] = 8'h6c;
            8'hb : a[0:7] = 8'h62;
            8'hc : a[0:7] = 8'h48;
            8'hd : a[0:7] = 8'h46;
            8'he : a[0:7] = 8'h54;
            8'hf : a[0:7] = 8'h5a;
            8'h10 : a[0:7] = 8'he0;
            8'h11 : a[0:7] = 8'hee;
            8'h12 : a[0:7] = 8'hfc;
            8'h13 : a[0:7] = 8'hf2;
            8'h14 : a[0:7] = 8'hd8;
            8'h15 : a[0:7] = 8'hd6;
            8'h16 : a[0:7] = 8'hc4;
            8'h17 : a[0:7] = 8'hca;
            8'h18 : a[0:7] = 8'h90;
            8'h19 : a[0:7] = 8'h9e;
            8'h1a : a[0:7] = 8'h8c;
            8'h1b : a[0:7] = 8'h82;
            8'h1c : a[0:7] = 8'ha8;
            8'h1d : a[0:7] = 8'ha6;
            8'h1e : a[0:7] = 8'hb4;
            8'h1f : a[0:7] = 8'hba;
            8'h20 : a[0:7] = 8'hdb;
            8'h21 : a[0:7] = 8'hd5;
            8'h22 : a[0:7] = 8'hc7;
            8'h23 : a[0:7] = 8'hc9;
            8'h24 : a[0:7] = 8'he3;
            8'h25 : a[0:7] = 8'hed;
            8'h26 : a[0:7] = 8'hff;
            8'h27 : a[0:7] = 8'hf1;
            8'h28 : a[0:7] = 8'hab;
            8'h29 : a[0:7] = 8'ha5;
            8'h2a : a[0:7] = 8'hb7;
            8'h2b : a[0:7] = 8'hb9;
            8'h2c : a[0:7] = 8'h93;
            8'h2d : a[0:7] = 8'h9d;
            8'h2e : a[0:7] = 8'h8f;
            8'h2f : a[0:7] = 8'h81;
            8'h30 : a[0:7] = 8'h3b;
            8'h31 : a[0:7] = 8'h35;
            8'h32 : a[0:7] = 8'h27;
            8'h33 : a[0:7] = 8'h29;
            8'h34 : a[0:7] = 8'h3;
            8'h35 : a[0:7] = 8'hd;
            8'h36 : a[0:7] = 8'h1f;
            8'h37 : a[0:7] = 8'h11;
            8'h38 : a[0:7] = 8'h4b;
            8'h39 : a[0:7] = 8'h45;
            8'h3a : a[0:7] = 8'h57;
            8'h3b : a[0:7] = 8'h59;
            8'h3c : a[0:7] = 8'h73;
            8'h3d : a[0:7] = 8'h7d;
            8'h3e : a[0:7] = 8'h6f;
            8'h3f : a[0:7] = 8'h61;
            8'h40 : a[0:7] = 8'had;
            8'h41 : a[0:7] = 8'ha3;
            8'h42 : a[0:7] = 8'hb1;
            8'h43 : a[0:7] = 8'hbf;
            8'h44 : a[0:7] = 8'h95;
            8'h45 : a[0:7] = 8'h9b;
            8'h46 : a[0:7] = 8'h89;
            8'h47 : a[0:7] = 8'h87;
            8'h48 : a[0:7] = 8'hdd;
            8'h49 : a[0:7] = 8'hd3;
            8'h4a : a[0:7] = 8'hc1;
            8'h4b : a[0:7] = 8'hcf;
            8'h4c : a[0:7] = 8'he5;
            8'h4d : a[0:7] = 8'heb;
            8'h4e : a[0:7] = 8'hf9;
            8'h4f : a[0:7] = 8'hf7;
            8'h50 : a[0:7] = 8'h4d;
            8'h51 : a[0:7] = 8'h43;
            8'h52 : a[0:7] = 8'h51;
            8'h53 : a[0:7] = 8'h5f;
            8'h54 : a[0:7] = 8'h75;
            8'h55 : a[0:7] = 8'h7b;
            8'h56 : a[0:7] = 8'h69;
            8'h57 : a[0:7] = 8'h67;
            8'h58 : a[0:7] = 8'h3d;
            8'h59 : a[0:7] = 8'h33;
            8'h5a : a[0:7] = 8'h21;
            8'h5b : a[0:7] = 8'h2f;
            8'h5c : a[0:7] = 8'h5;
            8'h5d : a[0:7] = 8'hb;
            8'h5e : a[0:7] = 8'h19;
            8'h5f : a[0:7] = 8'h17;
            8'h60 : a[0:7] = 8'h76;
            8'h61 : a[0:7] = 8'h78;
            8'h62 : a[0:7] = 8'h6a;
            8'h63 : a[0:7] = 8'h64;
            8'h64 : a[0:7] = 8'h4e;
            8'h65 : a[0:7] = 8'h40;
            8'h66 : a[0:7] = 8'h52;
            8'h67 : a[0:7] = 8'h5c;
            8'h68 : a[0:7] = 8'h6;
            8'h69 : a[0:7] = 8'h8;
            8'h6a : a[0:7] = 8'h1a;
            8'h6b : a[0:7] = 8'h14;
            8'h6c : a[0:7] = 8'h3e;
            8'h6d : a[0:7] = 8'h30;
            8'h6e : a[0:7] = 8'h22;
            8'h6f : a[0:7] = 8'h2c;
            8'h70 : a[0:7] = 8'h96;
            8'h71 : a[0:7] = 8'h98;
            8'h72 : a[0:7] = 8'h8a;
            8'h73 : a[0:7] = 8'h84;
            8'h74 : a[0:7] = 8'hae;
            8'h75 : a[0:7] = 8'ha0;
            8'h76 : a[0:7] = 8'hb2;
            8'h77 : a[0:7] = 8'hbc;
            8'h78 : a[0:7] = 8'he6;
            8'h79 : a[0:7] = 8'he8;
            8'h7a : a[0:7] = 8'hfa;
            8'h7b : a[0:7] = 8'hf4;
            8'h7c : a[0:7] = 8'hde;
            8'h7d : a[0:7] = 8'hd0;
            8'h7e : a[0:7] = 8'hc2;
            8'h7f : a[0:7] = 8'hcc;
            8'h80 : a[0:7] = 8'h41;
            8'h81 : a[0:7] = 8'h4f;
            8'h82 : a[0:7] = 8'h5d;
            8'h83 : a[0:7] = 8'h53;
            8'h84 : a[0:7] = 8'h79;
            8'h85 : a[0:7] = 8'h77;
            8'h86 : a[0:7] = 8'h65;
            8'h87 : a[0:7] = 8'h6b;
            8'h88 : a[0:7] = 8'h31;
            8'h89 : a[0:7] = 8'h3f;
            8'h8a : a[0:7] = 8'h2d;
            8'h8b : a[0:7] = 8'h23;
            8'h8c : a[0:7] = 8'h9;
            8'h8d : a[0:7] = 8'h7;
            8'h8e : a[0:7] = 8'h15;
            8'h8f : a[0:7] = 8'h1b;
            8'h90 : a[0:7] = 8'ha1;
            8'h91 : a[0:7] = 8'haf;
            8'h92 : a[0:7] = 8'hbd;
            8'h93 : a[0:7] = 8'hb3;
            8'h94 : a[0:7] = 8'h99;
            8'h95 : a[0:7] = 8'h97;
            8'h96 : a[0:7] = 8'h85;
            8'h97 : a[0:7] = 8'h8b;
            8'h98 : a[0:7] = 8'hd1;
            8'h99 : a[0:7] = 8'hdf;
            8'h9a : a[0:7] = 8'hcd;
            8'h9b : a[0:7] = 8'hc3;
            8'h9c : a[0:7] = 8'he9;
            8'h9d : a[0:7] = 8'he7;
            8'h9e : a[0:7] = 8'hf5;
            8'h9f : a[0:7] = 8'hfb;
            8'ha0 : a[0:7] = 8'h9a;
            8'ha1 : a[0:7] = 8'h94;
            8'ha2 : a[0:7] = 8'h86;
            8'ha3 : a[0:7] = 8'h88;
            8'ha4 : a[0:7] = 8'ha2;
            8'ha5 : a[0:7] = 8'hac;
            8'ha6 : a[0:7] = 8'hbe;
            8'ha7 : a[0:7] = 8'hb0;
            8'ha8 : a[0:7] = 8'hea;
            8'ha9 : a[0:7] = 8'he4;
            8'haa : a[0:7] = 8'hf6;
            8'hab : a[0:7] = 8'hf8;
            8'hac : a[0:7] = 8'hd2;
            8'had : a[0:7] = 8'hdc;
            8'hae : a[0:7] = 8'hce;
            8'haf : a[0:7] = 8'hc0;
            8'hb0 : a[0:7] = 8'h7a;
            8'hb1 : a[0:7] = 8'h74;
            8'hb2 : a[0:7] = 8'h66;
            8'hb3 : a[0:7] = 8'h68;
            8'hb4 : a[0:7] = 8'h42;
            8'hb5 : a[0:7] = 8'h4c;
            8'hb6 : a[0:7] = 8'h5e;
            8'hb7 : a[0:7] = 8'h50;
            8'hb8 : a[0:7] = 8'ha;
            8'hb9 : a[0:7] = 8'h4;
            8'hba : a[0:7] = 8'h16;
            8'hbb : a[0:7] = 8'h18;
            8'hbc : a[0:7] = 8'h32;
            8'hbd : a[0:7] = 8'h3c;
            8'hbe : a[0:7] = 8'h2e;
            8'hbf : a[0:7] = 8'h20;
            8'hc0 : a[0:7] = 8'hec;
            8'hc1 : a[0:7] = 8'he2;
            8'hc2 : a[0:7] = 8'hf0;
            8'hc3 : a[0:7] = 8'hfe;
            8'hc4 : a[0:7] = 8'hd4;
            8'hc5 : a[0:7] = 8'hda;
            8'hc6 : a[0:7] = 8'hc8;
            8'hc7 : a[0:7] = 8'hc6;
            8'hc8 : a[0:7] = 8'h9c;
            8'hc9 : a[0:7] = 8'h92;
            8'hca : a[0:7] = 8'h80;
            8'hcb : a[0:7] = 8'h8e;
            8'hcc : a[0:7] = 8'ha4;
            8'hcd : a[0:7] = 8'haa;
            8'hce : a[0:7] = 8'hb8;
            8'hcf : a[0:7] = 8'hb6;
            8'hd0 : a[0:7] = 8'hc;
            8'hd1 : a[0:7] = 8'h2;
            8'hd2 : a[0:7] = 8'h10;
            8'hd3 : a[0:7] = 8'h1e;
            8'hd4 : a[0:7] = 8'h34;
            8'hd5 : a[0:7] = 8'h3a;
            8'hd6 : a[0:7] = 8'h28;
            8'hd7 : a[0:7] = 8'h26;
            8'hd8 : a[0:7] = 8'h7c;
            8'hd9 : a[0:7] = 8'h72;
            8'hda : a[0:7] = 8'h60;
            8'hdb : a[0:7] = 8'h6e;
            8'hdc : a[0:7] = 8'h44;
            8'hdd : a[0:7] = 8'h4a;
            8'hde : a[0:7] = 8'h58;
            8'hdf : a[0:7] = 8'h56;
            8'he0 : a[0:7] = 8'h37;
            8'he1 : a[0:7] = 8'h39;
            8'he2 : a[0:7] = 8'h2b;
            8'he3 : a[0:7] = 8'h25;
            8'he4 : a[0:7] = 8'hf;
            8'he5 : a[0:7] = 8'h1;
            8'he6 : a[0:7] = 8'h13;
            8'he7 : a[0:7] = 8'h1d;
            8'he8 : a[0:7] = 8'h47;
            8'he9 : a[0:7] = 8'h49;
            8'hea : a[0:7] = 8'h5b;
            8'heb : a[0:7] = 8'h55;
            8'hec : a[0:7] = 8'h7f;
            8'hed : a[0:7] = 8'h71;
            8'hee : a[0:7] = 8'h63;
            8'hef : a[0:7] = 8'h6d;
            8'hf0 : a[0:7] = 8'hd7;
            8'hf1 : a[0:7] = 8'hd9;
            8'hf2 : a[0:7] = 8'hcb;
            8'hf3 : a[0:7] = 8'hc5;
            8'hf4 : a[0:7] = 8'hef;
            8'hf5 : a[0:7] = 8'he1;
            8'hf6 : a[0:7] = 8'hf3;
            8'hf7 : a[0:7] = 8'hfd;
            8'hf8 : a[0:7] = 8'ha7;
            8'hf9 : a[0:7] = 8'ha9;
            8'hfa : a[0:7] = 8'hbb;
            8'hfb : a[0:7] = 8'hb5;
            8'hfc : a[0:7] = 8'h9f;
            8'hfd : a[0:7] = 8'h91;
            8'hfe : a[0:7] = 8'h83;
            8'hff : a[0:7] = 8'h8d;
        endcase
    end

    // Multiplication with 11
    always @(row[8:15]) begin
        case (row[8:15])
            8'h0 : b[0:7] = 8'h0;
            8'h1 : b[0:7] = 8'hb;
            8'h2 : b[0:7] = 8'h16;
            8'h3 : b[0:7] = 8'h1d;
            8'h4 : b[0:7] = 8'h2c;
            8'h5 : b[0:7] = 8'h27;
            8'h6 : b[0:7] = 8'h3a;
            8'h7 : b[0:7] = 8'h31;
            8'h8 : b[0:7] = 8'h58;
            8'h9 : b[0:7] = 8'h53;
            8'ha : b[0:7] = 8'h4e;
            8'hb : b[0:7] = 8'h45;
            8'hc : b[0:7] = 8'h74;
            8'hd : b[0:7] = 8'h7f;
            8'he : b[0:7] = 8'h62;
            8'hf : b[0:7] = 8'h69;
            8'h10 : b[0:7] = 8'hb0;
            8'h11 : b[0:7] = 8'hbb;
            8'h12 : b[0:7] = 8'ha6;
            8'h13 : b[0:7] = 8'had;
            8'h14 : b[0:7] = 8'h9c;
            8'h15 : b[0:7] = 8'h97;
            8'h16 : b[0:7] = 8'h8a;
            8'h17 : b[0:7] = 8'h81;
            8'h18 : b[0:7] = 8'he8;
            8'h19 : b[0:7] = 8'he3;
            8'h1a : b[0:7] = 8'hfe;
            8'h1b : b[0:7] = 8'hf5;
            8'h1c : b[0:7] = 8'hc4;
            8'h1d : b[0:7] = 8'hcf;
            8'h1e : b[0:7] = 8'hd2;
            8'h1f : b[0:7] = 8'hd9;
            8'h20 : b[0:7] = 8'h7b;
            8'h21 : b[0:7] = 8'h70;
            8'h22 : b[0:7] = 8'h6d;
            8'h23 : b[0:7] = 8'h66;
            8'h24 : b[0:7] = 8'h57;
            8'h25 : b[0:7] = 8'h5c;
            8'h26 : b[0:7] = 8'h41;
            8'h27 : b[0:7] = 8'h4a;
            8'h28 : b[0:7] = 8'h23;
            8'h29 : b[0:7] = 8'h28;
            8'h2a : b[0:7] = 8'h35;
            8'h2b : b[0:7] = 8'h3e;
            8'h2c : b[0:7] = 8'hf;
            8'h2d : b[0:7] = 8'h4;
            8'h2e : b[0:7] = 8'h19;
            8'h2f : b[0:7] = 8'h12;
            8'h30 : b[0:7] = 8'hcb;
            8'h31 : b[0:7] = 8'hc0;
            8'h32 : b[0:7] = 8'hdd;
            8'h33 : b[0:7] = 8'hd6;
            8'h34 : b[0:7] = 8'he7;
            8'h35 : b[0:7] = 8'hec;
            8'h36 : b[0:7] = 8'hf1;
            8'h37 : b[0:7] = 8'hfa;
            8'h38 : b[0:7] = 8'h93;
            8'h39 : b[0:7] = 8'h98;
            8'h3a : b[0:7] = 8'h85;
            8'h3b : b[0:7] = 8'h8e;
            8'h3c : b[0:7] = 8'hbf;
            8'h3d : b[0:7] = 8'hb4;
            8'h3e : b[0:7] = 8'ha9;
            8'h3f : b[0:7] = 8'ha2;
            8'h40 : b[0:7] = 8'hf6;
            8'h41 : b[0:7] = 8'hfd;
            8'h42 : b[0:7] = 8'he0;
            8'h43 : b[0:7] = 8'heb;
            8'h44 : b[0:7] = 8'hda;
            8'h45 : b[0:7] = 8'hd1;
            8'h46 : b[0:7] = 8'hcc;
            8'h47 : b[0:7] = 8'hc7;
            8'h48 : b[0:7] = 8'hae;
            8'h49 : b[0:7] = 8'ha5;
            8'h4a : b[0:7] = 8'hb8;
            8'h4b : b[0:7] = 8'hb3;
            8'h4c : b[0:7] = 8'h82;
            8'h4d : b[0:7] = 8'h89;
            8'h4e : b[0:7] = 8'h94;
            8'h4f : b[0:7] = 8'h9f;
            8'h50 : b[0:7] = 8'h46;
            8'h51 : b[0:7] = 8'h4d;
            8'h52 : b[0:7] = 8'h50;
            8'h53 : b[0:7] = 8'h5b;
            8'h54 : b[0:7] = 8'h6a;
            8'h55 : b[0:7] = 8'h61;
            8'h56 : b[0:7] = 8'h7c;
            8'h57 : b[0:7] = 8'h77;
            8'h58 : b[0:7] = 8'h1e;
            8'h59 : b[0:7] = 8'h15;
            8'h5a : b[0:7] = 8'h8;
            8'h5b : b[0:7] = 8'h3;
            8'h5c : b[0:7] = 8'h32;
            8'h5d : b[0:7] = 8'h39;
            8'h5e : b[0:7] = 8'h24;
            8'h5f : b[0:7] = 8'h2f;
            8'h60 : b[0:7] = 8'h8d;
            8'h61 : b[0:7] = 8'h86;
            8'h62 : b[0:7] = 8'h9b;
            8'h63 : b[0:7] = 8'h90;
            8'h64 : b[0:7] = 8'ha1;
            8'h65 : b[0:7] = 8'haa;
            8'h66 : b[0:7] = 8'hb7;
            8'h67 : b[0:7] = 8'hbc;
            8'h68 : b[0:7] = 8'hd5;
            8'h69 : b[0:7] = 8'hde;
            8'h6a : b[0:7] = 8'hc3;
            8'h6b : b[0:7] = 8'hc8;
            8'h6c : b[0:7] = 8'hf9;
            8'h6d : b[0:7] = 8'hf2;
            8'h6e : b[0:7] = 8'hef;
            8'h6f : b[0:7] = 8'he4;
            8'h70 : b[0:7] = 8'h3d;
            8'h71 : b[0:7] = 8'h36;
            8'h72 : b[0:7] = 8'h2b;
            8'h73 : b[0:7] = 8'h20;
            8'h74 : b[0:7] = 8'h11;
            8'h75 : b[0:7] = 8'h1a;
            8'h76 : b[0:7] = 8'h7;
            8'h77 : b[0:7] = 8'hc;
            8'h78 : b[0:7] = 8'h65;
            8'h79 : b[0:7] = 8'h6e;
            8'h7a : b[0:7] = 8'h73;
            8'h7b : b[0:7] = 8'h78;
            8'h7c : b[0:7] = 8'h49;
            8'h7d : b[0:7] = 8'h42;
            8'h7e : b[0:7] = 8'h5f;
            8'h7f : b[0:7] = 8'h54;
            8'h80 : b[0:7] = 8'hf7;
            8'h81 : b[0:7] = 8'hfc;
            8'h82 : b[0:7] = 8'he1;
            8'h83 : b[0:7] = 8'hea;
            8'h84 : b[0:7] = 8'hdb;
            8'h85 : b[0:7] = 8'hd0;
            8'h86 : b[0:7] = 8'hcd;
            8'h87 : b[0:7] = 8'hc6;
            8'h88 : b[0:7] = 8'haf;
            8'h89 : b[0:7] = 8'ha4;
            8'h8a : b[0:7] = 8'hb9;
            8'h8b : b[0:7] = 8'hb2;
            8'h8c : b[0:7] = 8'h83;
            8'h8d : b[0:7] = 8'h88;
            8'h8e : b[0:7] = 8'h95;
            8'h8f : b[0:7] = 8'h9e;
            8'h90 : b[0:7] = 8'h47;
            8'h91 : b[0:7] = 8'h4c;
            8'h92 : b[0:7] = 8'h51;
            8'h93 : b[0:7] = 8'h5a;
            8'h94 : b[0:7] = 8'h6b;
            8'h95 : b[0:7] = 8'h60;
            8'h96 : b[0:7] = 8'h7d;
            8'h97 : b[0:7] = 8'h76;
            8'h98 : b[0:7] = 8'h1f;
            8'h99 : b[0:7] = 8'h14;
            8'h9a : b[0:7] = 8'h9;
            8'h9b : b[0:7] = 8'h2;
            8'h9c : b[0:7] = 8'h33;
            8'h9d : b[0:7] = 8'h38;
            8'h9e : b[0:7] = 8'h25;
            8'h9f : b[0:7] = 8'h2e;
            8'ha0 : b[0:7] = 8'h8c;
            8'ha1 : b[0:7] = 8'h87;
            8'ha2 : b[0:7] = 8'h9a;
            8'ha3 : b[0:7] = 8'h91;
            8'ha4 : b[0:7] = 8'ha0;
            8'ha5 : b[0:7] = 8'hab;
            8'ha6 : b[0:7] = 8'hb6;
            8'ha7 : b[0:7] = 8'hbd;
            8'ha8 : b[0:7] = 8'hd4;
            8'ha9 : b[0:7] = 8'hdf;
            8'haa : b[0:7] = 8'hc2;
            8'hab : b[0:7] = 8'hc9;
            8'hac : b[0:7] = 8'hf8;
            8'had : b[0:7] = 8'hf3;
            8'hae : b[0:7] = 8'hee;
            8'haf : b[0:7] = 8'he5;
            8'hb0 : b[0:7] = 8'h3c;
            8'hb1 : b[0:7] = 8'h37;
            8'hb2 : b[0:7] = 8'h2a;
            8'hb3 : b[0:7] = 8'h21;
            8'hb4 : b[0:7] = 8'h10;
            8'hb5 : b[0:7] = 8'h1b;
            8'hb6 : b[0:7] = 8'h6;
            8'hb7 : b[0:7] = 8'hd;
            8'hb8 : b[0:7] = 8'h64;
            8'hb9 : b[0:7] = 8'h6f;
            8'hba : b[0:7] = 8'h72;
            8'hbb : b[0:7] = 8'h79;
            8'hbc : b[0:7] = 8'h48;
            8'hbd : b[0:7] = 8'h43;
            8'hbe : b[0:7] = 8'h5e;
            8'hbf : b[0:7] = 8'h55;
            8'hc0 : b[0:7] = 8'h1;
            8'hc1 : b[0:7] = 8'ha;
            8'hc2 : b[0:7] = 8'h17;
            8'hc3 : b[0:7] = 8'h1c;
            8'hc4 : b[0:7] = 8'h2d;
            8'hc5 : b[0:7] = 8'h26;
            8'hc6 : b[0:7] = 8'h3b;
            8'hc7 : b[0:7] = 8'h30;
            8'hc8 : b[0:7] = 8'h59;
            8'hc9 : b[0:7] = 8'h52;
            8'hca : b[0:7] = 8'h4f;
            8'hcb : b[0:7] = 8'h44;
            8'hcc : b[0:7] = 8'h75;
            8'hcd : b[0:7] = 8'h7e;
            8'hce : b[0:7] = 8'h63;
            8'hcf : b[0:7] = 8'h68;
            8'hd0 : b[0:7] = 8'hb1;
            8'hd1 : b[0:7] = 8'hba;
            8'hd2 : b[0:7] = 8'ha7;
            8'hd3 : b[0:7] = 8'hac;
            8'hd4 : b[0:7] = 8'h9d;
            8'hd5 : b[0:7] = 8'h96;
            8'hd6 : b[0:7] = 8'h8b;
            8'hd7 : b[0:7] = 8'h80;
            8'hd8 : b[0:7] = 8'he9;
            8'hd9 : b[0:7] = 8'he2;
            8'hda : b[0:7] = 8'hff;
            8'hdb : b[0:7] = 8'hf4;
            8'hdc : b[0:7] = 8'hc5;
            8'hdd : b[0:7] = 8'hce;
            8'hde : b[0:7] = 8'hd3;
            8'hdf : b[0:7] = 8'hd8;
            8'he0 : b[0:7] = 8'h7a;
            8'he1 : b[0:7] = 8'h71;
            8'he2 : b[0:7] = 8'h6c;
            8'he3 : b[0:7] = 8'h67;
            8'he4 : b[0:7] = 8'h56;
            8'he5 : b[0:7] = 8'h5d;
            8'he6 : b[0:7] = 8'h40;
            8'he7 : b[0:7] = 8'h4b;
            8'he8 : b[0:7] = 8'h22;
            8'he9 : b[0:7] = 8'h29;
            8'hea : b[0:7] = 8'h34;
            8'heb : b[0:7] = 8'h3f;
            8'hec : b[0:7] = 8'he;
            8'hed : b[0:7] = 8'h5;
            8'hee : b[0:7] = 8'h18;
            8'hef : b[0:7] = 8'h13;
            8'hf0 : b[0:7] = 8'hca;
            8'hf1 : b[0:7] = 8'hc1;
            8'hf2 : b[0:7] = 8'hdc;
            8'hf3 : b[0:7] = 8'hd7;
            8'hf4 : b[0:7] = 8'he6;
            8'hf5 : b[0:7] = 8'hed;
            8'hf6 : b[0:7] = 8'hf0;
            8'hf7 : b[0:7] = 8'hfb;
            8'hf8 : b[0:7] = 8'h92;
            8'hf9 : b[0:7] = 8'h99;
            8'hfa : b[0:7] = 8'h84;
            8'hfb : b[0:7] = 8'h8f;
            8'hfc : b[0:7] = 8'hbe;
            8'hfd : b[0:7] = 8'hb5;
            8'hfe : b[0:7] = 8'ha8;
            8'hff : b[0:7] = 8'ha3;
        endcase
    end

    // Multiplication with 13
    always @(row[16:23]) begin
        case (row[16:23])
			8'h0 : c[0:7] = 8'h0;
			8'h1 : c[0:7] = 8'hd;
			8'h2 : c[0:7] = 8'h1a;
			8'h3 : c[0:7] = 8'h17;
			8'h4 : c[0:7] = 8'h34;
			8'h5 : c[0:7] = 8'h39;
			8'h6 : c[0:7] = 8'h2e;
			8'h7 : c[0:7] = 8'h23;
			8'h8 : c[0:7] = 8'h68;
			8'h9 : c[0:7] = 8'h65;
			8'ha : c[0:7] = 8'h72;
			8'hb : c[0:7] = 8'h7f;
			8'hc : c[0:7] = 8'h5c;
			8'hd : c[0:7] = 8'h51;
			8'he : c[0:7] = 8'h46;
			8'hf : c[0:7] = 8'h4b;
			8'h10 : c[0:7] = 8'hd0;
			8'h11 : c[0:7] = 8'hdd;
			8'h12 : c[0:7] = 8'hca;
			8'h13 : c[0:7] = 8'hc7;
			8'h14 : c[0:7] = 8'he4;
			8'h15 : c[0:7] = 8'he9;
			8'h16 : c[0:7] = 8'hfe;
			8'h17 : c[0:7] = 8'hf3;
			8'h18 : c[0:7] = 8'hb8;
			8'h19 : c[0:7] = 8'hb5;
			8'h1a : c[0:7] = 8'ha2;
			8'h1b : c[0:7] = 8'haf;
			8'h1c : c[0:7] = 8'h8c;
			8'h1d : c[0:7] = 8'h81;
			8'h1e : c[0:7] = 8'h96;
			8'h1f : c[0:7] = 8'h9b;
			8'h20 : c[0:7] = 8'hbb;
			8'h21 : c[0:7] = 8'hb6;
			8'h22 : c[0:7] = 8'ha1;
			8'h23 : c[0:7] = 8'hac;
			8'h24 : c[0:7] = 8'h8f;
			8'h25 : c[0:7] = 8'h82;
			8'h26 : c[0:7] = 8'h95;
			8'h27 : c[0:7] = 8'h98;
			8'h28 : c[0:7] = 8'hd3;
			8'h29 : c[0:7] = 8'hde;
			8'h2a : c[0:7] = 8'hc9;
			8'h2b : c[0:7] = 8'hc4;
			8'h2c : c[0:7] = 8'he7;
			8'h2d : c[0:7] = 8'hea;
			8'h2e : c[0:7] = 8'hfd;
			8'h2f : c[0:7] = 8'hf0;
			8'h30 : c[0:7] = 8'h6b;
			8'h31 : c[0:7] = 8'h66;
			8'h32 : c[0:7] = 8'h71;
			8'h33 : c[0:7] = 8'h7c;
			8'h34 : c[0:7] = 8'h5f;
			8'h35 : c[0:7] = 8'h52;
			8'h36 : c[0:7] = 8'h45;
			8'h37 : c[0:7] = 8'h48;
			8'h38 : c[0:7] = 8'h3;
			8'h39 : c[0:7] = 8'he;
			8'h3a : c[0:7] = 8'h19;
			8'h3b : c[0:7] = 8'h14;
			8'h3c : c[0:7] = 8'h37;
			8'h3d : c[0:7] = 8'h3a;
			8'h3e : c[0:7] = 8'h2d;
			8'h3f : c[0:7] = 8'h20;
			8'h40 : c[0:7] = 8'h6d;
			8'h41 : c[0:7] = 8'h60;
			8'h42 : c[0:7] = 8'h77;
			8'h43 : c[0:7] = 8'h7a;
			8'h44 : c[0:7] = 8'h59;
			8'h45 : c[0:7] = 8'h54;
			8'h46 : c[0:7] = 8'h43;
			8'h47 : c[0:7] = 8'h4e;
			8'h48 : c[0:7] = 8'h5;
			8'h49 : c[0:7] = 8'h8;
			8'h4a : c[0:7] = 8'h1f;
			8'h4b : c[0:7] = 8'h12;
			8'h4c : c[0:7] = 8'h31;
			8'h4d : c[0:7] = 8'h3c;
			8'h4e : c[0:7] = 8'h2b;
			8'h4f : c[0:7] = 8'h26;
			8'h50 : c[0:7] = 8'hbd;
			8'h51 : c[0:7] = 8'hb0;
			8'h52 : c[0:7] = 8'ha7;
			8'h53 : c[0:7] = 8'haa;
			8'h54 : c[0:7] = 8'h89;
			8'h55 : c[0:7] = 8'h84;
			8'h56 : c[0:7] = 8'h93;
			8'h57 : c[0:7] = 8'h9e;
			8'h58 : c[0:7] = 8'hd5;
			8'h59 : c[0:7] = 8'hd8;
			8'h5a : c[0:7] = 8'hcf;
			8'h5b : c[0:7] = 8'hc2;
			8'h5c : c[0:7] = 8'he1;
			8'h5d : c[0:7] = 8'hec;
			8'h5e : c[0:7] = 8'hfb;
			8'h5f : c[0:7] = 8'hf6;
			8'h60 : c[0:7] = 8'hd6;
			8'h61 : c[0:7] = 8'hdb;
			8'h62 : c[0:7] = 8'hcc;
			8'h63 : c[0:7] = 8'hc1;
			8'h64 : c[0:7] = 8'he2;
			8'h65 : c[0:7] = 8'hef;
			8'h66 : c[0:7] = 8'hf8;
			8'h67 : c[0:7] = 8'hf5;
			8'h68 : c[0:7] = 8'hbe;
			8'h69 : c[0:7] = 8'hb3;
			8'h6a : c[0:7] = 8'ha4;
			8'h6b : c[0:7] = 8'ha9;
			8'h6c : c[0:7] = 8'h8a;
			8'h6d : c[0:7] = 8'h87;
			8'h6e : c[0:7] = 8'h90;
			8'h6f : c[0:7] = 8'h9d;
			8'h70 : c[0:7] = 8'h6;
			8'h71 : c[0:7] = 8'hb;
			8'h72 : c[0:7] = 8'h1c;
			8'h73 : c[0:7] = 8'h11;
			8'h74 : c[0:7] = 8'h32;
			8'h75 : c[0:7] = 8'h3f;
			8'h76 : c[0:7] = 8'h28;
			8'h77 : c[0:7] = 8'h25;
			8'h78 : c[0:7] = 8'h6e;
			8'h79 : c[0:7] = 8'h63;
			8'h7a : c[0:7] = 8'h74;
			8'h7b : c[0:7] = 8'h79;
			8'h7c : c[0:7] = 8'h5a;
			8'h7d : c[0:7] = 8'h57;
			8'h7e : c[0:7] = 8'h40;
			8'h7f : c[0:7] = 8'h4d;
			8'h80 : c[0:7] = 8'hda;
			8'h81 : c[0:7] = 8'hd7;
			8'h82 : c[0:7] = 8'hc0;
			8'h83 : c[0:7] = 8'hcd;
			8'h84 : c[0:7] = 8'hee;
			8'h85 : c[0:7] = 8'he3;
			8'h86 : c[0:7] = 8'hf4;
			8'h87 : c[0:7] = 8'hf9;
			8'h88 : c[0:7] = 8'hb2;
			8'h89 : c[0:7] = 8'hbf;
			8'h8a : c[0:7] = 8'ha8;
			8'h8b : c[0:7] = 8'ha5;
			8'h8c : c[0:7] = 8'h86;
			8'h8d : c[0:7] = 8'h8b;
			8'h8e : c[0:7] = 8'h9c;
			8'h8f : c[0:7] = 8'h91;
			8'h90 : c[0:7] = 8'ha;
			8'h91 : c[0:7] = 8'h7;
			8'h92 : c[0:7] = 8'h10;
			8'h93 : c[0:7] = 8'h1d;
			8'h94 : c[0:7] = 8'h3e;
			8'h95 : c[0:7] = 8'h33;
			8'h96 : c[0:7] = 8'h24;
			8'h97 : c[0:7] = 8'h29;
			8'h98 : c[0:7] = 8'h62;
			8'h99 : c[0:7] = 8'h6f;
			8'h9a : c[0:7] = 8'h78;
			8'h9b : c[0:7] = 8'h75;
			8'h9c : c[0:7] = 8'h56;
			8'h9d : c[0:7] = 8'h5b;
			8'h9e : c[0:7] = 8'h4c;
			8'h9f : c[0:7] = 8'h41;
			8'ha0 : c[0:7] = 8'h61;
			8'ha1 : c[0:7] = 8'h6c;
			8'ha2 : c[0:7] = 8'h7b;
			8'ha3 : c[0:7] = 8'h76;
			8'ha4 : c[0:7] = 8'h55;
			8'ha5 : c[0:7] = 8'h58;
			8'ha6 : c[0:7] = 8'h4f;
			8'ha7 : c[0:7] = 8'h42;
			8'ha8 : c[0:7] = 8'h9;
			8'ha9 : c[0:7] = 8'h4;
			8'haa : c[0:7] = 8'h13;
			8'hab : c[0:7] = 8'h1e;
			8'hac : c[0:7] = 8'h3d;
			8'had : c[0:7] = 8'h30;
			8'hae : c[0:7] = 8'h27;
			8'haf : c[0:7] = 8'h2a;
			8'hb0 : c[0:7] = 8'hb1;
			8'hb1 : c[0:7] = 8'hbc;
			8'hb2 : c[0:7] = 8'hab;
			8'hb3 : c[0:7] = 8'ha6;
			8'hb4 : c[0:7] = 8'h85;
			8'hb5 : c[0:7] = 8'h88;
			8'hb6 : c[0:7] = 8'h9f;
			8'hb7 : c[0:7] = 8'h92;
			8'hb8 : c[0:7] = 8'hd9;
			8'hb9 : c[0:7] = 8'hd4;
			8'hba : c[0:7] = 8'hc3;
			8'hbb : c[0:7] = 8'hce;
			8'hbc : c[0:7] = 8'hed;
			8'hbd : c[0:7] = 8'he0;
			8'hbe : c[0:7] = 8'hf7;
			8'hbf : c[0:7] = 8'hfa;
			8'hc0 : c[0:7] = 8'hb7;
			8'hc1 : c[0:7] = 8'hba;
			8'hc2 : c[0:7] = 8'had;
			8'hc3 : c[0:7] = 8'ha0;
			8'hc4 : c[0:7] = 8'h83;
			8'hc5 : c[0:7] = 8'h8e;
			8'hc6 : c[0:7] = 8'h99;
			8'hc7 : c[0:7] = 8'h94;
			8'hc8 : c[0:7] = 8'hdf;
			8'hc9 : c[0:7] = 8'hd2;
			8'hca : c[0:7] = 8'hc5;
			8'hcb : c[0:7] = 8'hc8;
			8'hcc : c[0:7] = 8'heb;
			8'hcd : c[0:7] = 8'he6;
			8'hce : c[0:7] = 8'hf1;
			8'hcf : c[0:7] = 8'hfc;
			8'hd0 : c[0:7] = 8'h67;
			8'hd1 : c[0:7] = 8'h6a;
			8'hd2 : c[0:7] = 8'h7d;
			8'hd3 : c[0:7] = 8'h70;
			8'hd4 : c[0:7] = 8'h53;
			8'hd5 : c[0:7] = 8'h5e;
			8'hd6 : c[0:7] = 8'h49;
			8'hd7 : c[0:7] = 8'h44;
			8'hd8 : c[0:7] = 8'hf;
			8'hd9 : c[0:7] = 8'h2;
			8'hda : c[0:7] = 8'h15;
			8'hdb : c[0:7] = 8'h18;
			8'hdc : c[0:7] = 8'h3b;
			8'hdd : c[0:7] = 8'h36;
			8'hde : c[0:7] = 8'h21;
			8'hdf : c[0:7] = 8'h2c;
			8'he0 : c[0:7] = 8'hc;
			8'he1 : c[0:7] = 8'h1;
			8'he2 : c[0:7] = 8'h16;
			8'he3 : c[0:7] = 8'h1b;
			8'he4 : c[0:7] = 8'h38;
			8'he5 : c[0:7] = 8'h35;
			8'he6 : c[0:7] = 8'h22;
			8'he7 : c[0:7] = 8'h2f;
			8'he8 : c[0:7] = 8'h64;
			8'he9 : c[0:7] = 8'h69;
			8'hea : c[0:7] = 8'h7e;
			8'heb : c[0:7] = 8'h73;
			8'hec : c[0:7] = 8'h50;
			8'hed : c[0:7] = 8'h5d;
			8'hee : c[0:7] = 8'h4a;
			8'hef : c[0:7] = 8'h47;
			8'hf0 : c[0:7] = 8'hdc;
			8'hf1 : c[0:7] = 8'hd1;
			8'hf2 : c[0:7] = 8'hc6;
			8'hf3 : c[0:7] = 8'hcb;
			8'hf4 : c[0:7] = 8'he8;
			8'hf5 : c[0:7] = 8'he5;
			8'hf6 : c[0:7] = 8'hf2;
			8'hf7 : c[0:7] = 8'hff;
			8'hf8 : c[0:7] = 8'hb4;
			8'hf9 : c[0:7] = 8'hb9;
			8'hfa : c[0:7] = 8'hae;
			8'hfb : c[0:7] = 8'ha3;
			8'hfc : c[0:7] = 8'h80;
			8'hfd : c[0:7] = 8'h8d;
			8'hfe : c[0:7] = 8'h9a;
			8'hff : c[0:7] = 8'h97;
        endcase
    end

    // Multiplication with 9
    always @(row[24:31]) begin
        case (row[24:31])
			8'h0 : d[0:7] = 8'h0;
			8'h1 : d[0:7] = 8'h9;
			8'h2 : d[0:7] = 8'h12;
			8'h3 : d[0:7] = 8'h1b;
			8'h4 : d[0:7] = 8'h24;
			8'h5 : d[0:7] = 8'h2d;
			8'h6 : d[0:7] = 8'h36;
			8'h7 : d[0:7] = 8'h3f;
			8'h8 : d[0:7] = 8'h48;
			8'h9 : d[0:7] = 8'h41;
			8'ha : d[0:7] = 8'h5a;
			8'hb : d[0:7] = 8'h53;
			8'hc : d[0:7] = 8'h6c;
			8'hd : d[0:7] = 8'h65;
			8'he : d[0:7] = 8'h7e;
			8'hf : d[0:7] = 8'h77;
			8'h10 : d[0:7] = 8'h90;
			8'h11 : d[0:7] = 8'h99;
			8'h12 : d[0:7] = 8'h82;
			8'h13 : d[0:7] = 8'h8b;
			8'h14 : d[0:7] = 8'hb4;
			8'h15 : d[0:7] = 8'hbd;
			8'h16 : d[0:7] = 8'ha6;
			8'h17 : d[0:7] = 8'haf;
			8'h18 : d[0:7] = 8'hd8;
			8'h19 : d[0:7] = 8'hd1;
			8'h1a : d[0:7] = 8'hca;
			8'h1b : d[0:7] = 8'hc3;
			8'h1c : d[0:7] = 8'hfc;
			8'h1d : d[0:7] = 8'hf5;
			8'h1e : d[0:7] = 8'hee;
			8'h1f : d[0:7] = 8'he7;
			8'h20 : d[0:7] = 8'h3b;
			8'h21 : d[0:7] = 8'h32;
			8'h22 : d[0:7] = 8'h29;
			8'h23 : d[0:7] = 8'h20;
			8'h24 : d[0:7] = 8'h1f;
			8'h25 : d[0:7] = 8'h16;
			8'h26 : d[0:7] = 8'hd;
			8'h27 : d[0:7] = 8'h4;
			8'h28 : d[0:7] = 8'h73;
			8'h29 : d[0:7] = 8'h7a;
			8'h2a : d[0:7] = 8'h61;
			8'h2b : d[0:7] = 8'h68;
			8'h2c : d[0:7] = 8'h57;
			8'h2d : d[0:7] = 8'h5e;
			8'h2e : d[0:7] = 8'h45;
			8'h2f : d[0:7] = 8'h4c;
			8'h30 : d[0:7] = 8'hab;
			8'h31 : d[0:7] = 8'ha2;
			8'h32 : d[0:7] = 8'hb9;
			8'h33 : d[0:7] = 8'hb0;
			8'h34 : d[0:7] = 8'h8f;
			8'h35 : d[0:7] = 8'h86;
			8'h36 : d[0:7] = 8'h9d;
			8'h37 : d[0:7] = 8'h94;
			8'h38 : d[0:7] = 8'he3;
			8'h39 : d[0:7] = 8'hea;
			8'h3a : d[0:7] = 8'hf1;
			8'h3b : d[0:7] = 8'hf8;
			8'h3c : d[0:7] = 8'hc7;
			8'h3d : d[0:7] = 8'hce;
			8'h3e : d[0:7] = 8'hd5;
			8'h3f : d[0:7] = 8'hdc;
			8'h40 : d[0:7] = 8'h76;
			8'h41 : d[0:7] = 8'h7f;
			8'h42 : d[0:7] = 8'h64;
			8'h43 : d[0:7] = 8'h6d;
			8'h44 : d[0:7] = 8'h52;
			8'h45 : d[0:7] = 8'h5b;
			8'h46 : d[0:7] = 8'h40;
			8'h47 : d[0:7] = 8'h49;
			8'h48 : d[0:7] = 8'h3e;
			8'h49 : d[0:7] = 8'h37;
			8'h4a : d[0:7] = 8'h2c;
			8'h4b : d[0:7] = 8'h25;
			8'h4c : d[0:7] = 8'h1a;
			8'h4d : d[0:7] = 8'h13;
			8'h4e : d[0:7] = 8'h8;
			8'h4f : d[0:7] = 8'h1;
			8'h50 : d[0:7] = 8'he6;
			8'h51 : d[0:7] = 8'hef;
			8'h52 : d[0:7] = 8'hf4;
			8'h53 : d[0:7] = 8'hfd;
			8'h54 : d[0:7] = 8'hc2;
			8'h55 : d[0:7] = 8'hcb;
			8'h56 : d[0:7] = 8'hd0;
			8'h57 : d[0:7] = 8'hd9;
			8'h58 : d[0:7] = 8'hae;
			8'h59 : d[0:7] = 8'ha7;
			8'h5a : d[0:7] = 8'hbc;
			8'h5b : d[0:7] = 8'hb5;
			8'h5c : d[0:7] = 8'h8a;
			8'h5d : d[0:7] = 8'h83;
			8'h5e : d[0:7] = 8'h98;
			8'h5f : d[0:7] = 8'h91;
			8'h60 : d[0:7] = 8'h4d;
			8'h61 : d[0:7] = 8'h44;
			8'h62 : d[0:7] = 8'h5f;
			8'h63 : d[0:7] = 8'h56;
			8'h64 : d[0:7] = 8'h69;
			8'h65 : d[0:7] = 8'h60;
			8'h66 : d[0:7] = 8'h7b;
			8'h67 : d[0:7] = 8'h72;
			8'h68 : d[0:7] = 8'h5;
			8'h69 : d[0:7] = 8'hc;
			8'h6a : d[0:7] = 8'h17;
			8'h6b : d[0:7] = 8'h1e;
			8'h6c : d[0:7] = 8'h21;
			8'h6d : d[0:7] = 8'h28;
			8'h6e : d[0:7] = 8'h33;
			8'h6f : d[0:7] = 8'h3a;
			8'h70 : d[0:7] = 8'hdd;
			8'h71 : d[0:7] = 8'hd4;
			8'h72 : d[0:7] = 8'hcf;
			8'h73 : d[0:7] = 8'hc6;
			8'h74 : d[0:7] = 8'hf9;
			8'h75 : d[0:7] = 8'hf0;
			8'h76 : d[0:7] = 8'heb;
			8'h77 : d[0:7] = 8'he2;
			8'h78 : d[0:7] = 8'h95;
			8'h79 : d[0:7] = 8'h9c;
			8'h7a : d[0:7] = 8'h87;
			8'h7b : d[0:7] = 8'h8e;
			8'h7c : d[0:7] = 8'hb1;
			8'h7d : d[0:7] = 8'hb8;
			8'h7e : d[0:7] = 8'ha3;
			8'h7f : d[0:7] = 8'haa;
			8'h80 : d[0:7] = 8'hec;
			8'h81 : d[0:7] = 8'he5;
			8'h82 : d[0:7] = 8'hfe;
			8'h83 : d[0:7] = 8'hf7;
			8'h84 : d[0:7] = 8'hc8;
			8'h85 : d[0:7] = 8'hc1;
			8'h86 : d[0:7] = 8'hda;
			8'h87 : d[0:7] = 8'hd3;
			8'h88 : d[0:7] = 8'ha4;
			8'h89 : d[0:7] = 8'had;
			8'h8a : d[0:7] = 8'hb6;
			8'h8b : d[0:7] = 8'hbf;
			8'h8c : d[0:7] = 8'h80;
			8'h8d : d[0:7] = 8'h89;
			8'h8e : d[0:7] = 8'h92;
			8'h8f : d[0:7] = 8'h9b;
			8'h90 : d[0:7] = 8'h7c;
			8'h91 : d[0:7] = 8'h75;
			8'h92 : d[0:7] = 8'h6e;
			8'h93 : d[0:7] = 8'h67;
			8'h94 : d[0:7] = 8'h58;
			8'h95 : d[0:7] = 8'h51;
			8'h96 : d[0:7] = 8'h4a;
			8'h97 : d[0:7] = 8'h43;
			8'h98 : d[0:7] = 8'h34;
			8'h99 : d[0:7] = 8'h3d;
			8'h9a : d[0:7] = 8'h26;
			8'h9b : d[0:7] = 8'h2f;
			8'h9c : d[0:7] = 8'h10;
			8'h9d : d[0:7] = 8'h19;
			8'h9e : d[0:7] = 8'h2;
			8'h9f : d[0:7] = 8'hb;
			8'ha0 : d[0:7] = 8'hd7;
			8'ha1 : d[0:7] = 8'hde;
			8'ha2 : d[0:7] = 8'hc5;
			8'ha3 : d[0:7] = 8'hcc;
			8'ha4 : d[0:7] = 8'hf3;
			8'ha5 : d[0:7] = 8'hfa;
			8'ha6 : d[0:7] = 8'he1;
			8'ha7 : d[0:7] = 8'he8;
			8'ha8 : d[0:7] = 8'h9f;
			8'ha9 : d[0:7] = 8'h96;
			8'haa : d[0:7] = 8'h8d;
			8'hab : d[0:7] = 8'h84;
			8'hac : d[0:7] = 8'hbb;
			8'had : d[0:7] = 8'hb2;
			8'hae : d[0:7] = 8'ha9;
			8'haf : d[0:7] = 8'ha0;
			8'hb0 : d[0:7] = 8'h47;
			8'hb1 : d[0:7] = 8'h4e;
			8'hb2 : d[0:7] = 8'h55;
			8'hb3 : d[0:7] = 8'h5c;
			8'hb4 : d[0:7] = 8'h63;
			8'hb5 : d[0:7] = 8'h6a;
			8'hb6 : d[0:7] = 8'h71;
			8'hb7 : d[0:7] = 8'h78;
			8'hb8 : d[0:7] = 8'hf;
			8'hb9 : d[0:7] = 8'h6;
			8'hba : d[0:7] = 8'h1d;
			8'hbb : d[0:7] = 8'h14;
			8'hbc : d[0:7] = 8'h2b;
			8'hbd : d[0:7] = 8'h22;
			8'hbe : d[0:7] = 8'h39;
			8'hbf : d[0:7] = 8'h30;
			8'hc0 : d[0:7] = 8'h9a;
			8'hc1 : d[0:7] = 8'h93;
			8'hc2 : d[0:7] = 8'h88;
			8'hc3 : d[0:7] = 8'h81;
			8'hc4 : d[0:7] = 8'hbe;
			8'hc5 : d[0:7] = 8'hb7;
			8'hc6 : d[0:7] = 8'hac;
			8'hc7 : d[0:7] = 8'ha5;
			8'hc8 : d[0:7] = 8'hd2;
			8'hc9 : d[0:7] = 8'hdb;
			8'hca : d[0:7] = 8'hc0;
			8'hcb : d[0:7] = 8'hc9;
			8'hcc : d[0:7] = 8'hf6;
			8'hcd : d[0:7] = 8'hff;
			8'hce : d[0:7] = 8'he4;
			8'hcf : d[0:7] = 8'hed;
			8'hd0 : d[0:7] = 8'ha;
			8'hd1 : d[0:7] = 8'h3;
			8'hd2 : d[0:7] = 8'h18;
			8'hd3 : d[0:7] = 8'h11;
			8'hd4 : d[0:7] = 8'h2e;
			8'hd5 : d[0:7] = 8'h27;
			8'hd6 : d[0:7] = 8'h3c;
			8'hd7 : d[0:7] = 8'h35;
			8'hd8 : d[0:7] = 8'h42;
			8'hd9 : d[0:7] = 8'h4b;
			8'hda : d[0:7] = 8'h50;
			8'hdb : d[0:7] = 8'h59;
			8'hdc : d[0:7] = 8'h66;
			8'hdd : d[0:7] = 8'h6f;
			8'hde : d[0:7] = 8'h74;
			8'hdf : d[0:7] = 8'h7d;
			8'he0 : d[0:7] = 8'ha1;
			8'he1 : d[0:7] = 8'ha8;
			8'he2 : d[0:7] = 8'hb3;
			8'he3 : d[0:7] = 8'hba;
			8'he4 : d[0:7] = 8'h85;
			8'he5 : d[0:7] = 8'h8c;
			8'he6 : d[0:7] = 8'h97;
			8'he7 : d[0:7] = 8'h9e;
			8'he8 : d[0:7] = 8'he9;
			8'he9 : d[0:7] = 8'he0;
			8'hea : d[0:7] = 8'hfb;
			8'heb : d[0:7] = 8'hf2;
			8'hec : d[0:7] = 8'hcd;
			8'hed : d[0:7] = 8'hc4;
			8'hee : d[0:7] = 8'hdf;
			8'hef : d[0:7] = 8'hd6;
			8'hf0 : d[0:7] = 8'h31;
			8'hf1 : d[0:7] = 8'h38;
			8'hf2 : d[0:7] = 8'h23;
			8'hf3 : d[0:7] = 8'h2a;
			8'hf4 : d[0:7] = 8'h15;
			8'hf5 : d[0:7] = 8'h1c;
			8'hf6 : d[0:7] = 8'h7;
			8'hf7 : d[0:7] = 8'he;
			8'hf8 : d[0:7] = 8'h79;
			8'hf9 : d[0:7] = 8'h70;
			8'hfa : d[0:7] = 8'h6b;
			8'hfb : d[0:7] = 8'h62;
			8'hfc : d[0:7] = 8'h5d;
			8'hfd : d[0:7] = 8'h54;
			8'hfe : d[0:7] = 8'h4f;
			8'hff : d[0:7] = 8'h46;
        endcase
    end

    assign output_row = a ^ b ^ c ^ d;
    
endmodule


module MixColumn2RowInverse (
    input wire [0:31] row,
    output wire [0:7] output_row
);
    reg [0:7] a, b, c, d;

    // Multiplication with 9
    always @(row[0:7]) begin
        case (row[0:7])
            8'h0 : d[0:7] = 8'h0;
			8'h1 : d[0:7] = 8'h9;
			8'h2 : d[0:7] = 8'h12;
			8'h3 : d[0:7] = 8'h1b;
			8'h4 : d[0:7] = 8'h24;
			8'h5 : d[0:7] = 8'h2d;
			8'h6 : d[0:7] = 8'h36;
			8'h7 : d[0:7] = 8'h3f;
			8'h8 : d[0:7] = 8'h48;
			8'h9 : d[0:7] = 8'h41;
			8'ha : d[0:7] = 8'h5a;
			8'hb : d[0:7] = 8'h53;
			8'hc : d[0:7] = 8'h6c;
			8'hd : d[0:7] = 8'h65;
			8'he : d[0:7] = 8'h7e;
			8'hf : d[0:7] = 8'h77;
			8'h10 : d[0:7] = 8'h90;
			8'h11 : d[0:7] = 8'h99;
			8'h12 : d[0:7] = 8'h82;
			8'h13 : d[0:7] = 8'h8b;
			8'h14 : d[0:7] = 8'hb4;
			8'h15 : d[0:7] = 8'hbd;
			8'h16 : d[0:7] = 8'ha6;
			8'h17 : d[0:7] = 8'haf;
			8'h18 : d[0:7] = 8'hd8;
			8'h19 : d[0:7] = 8'hd1;
			8'h1a : d[0:7] = 8'hca;
			8'h1b : d[0:7] = 8'hc3;
			8'h1c : d[0:7] = 8'hfc;
			8'h1d : d[0:7] = 8'hf5;
			8'h1e : d[0:7] = 8'hee;
			8'h1f : d[0:7] = 8'he7;
			8'h20 : d[0:7] = 8'h3b;
			8'h21 : d[0:7] = 8'h32;
			8'h22 : d[0:7] = 8'h29;
			8'h23 : d[0:7] = 8'h20;
			8'h24 : d[0:7] = 8'h1f;
			8'h25 : d[0:7] = 8'h16;
			8'h26 : d[0:7] = 8'hd;
			8'h27 : d[0:7] = 8'h4;
			8'h28 : d[0:7] = 8'h73;
			8'h29 : d[0:7] = 8'h7a;
			8'h2a : d[0:7] = 8'h61;
			8'h2b : d[0:7] = 8'h68;
			8'h2c : d[0:7] = 8'h57;
			8'h2d : d[0:7] = 8'h5e;
			8'h2e : d[0:7] = 8'h45;
			8'h2f : d[0:7] = 8'h4c;
			8'h30 : d[0:7] = 8'hab;
			8'h31 : d[0:7] = 8'ha2;
			8'h32 : d[0:7] = 8'hb9;
			8'h33 : d[0:7] = 8'hb0;
			8'h34 : d[0:7] = 8'h8f;
			8'h35 : d[0:7] = 8'h86;
			8'h36 : d[0:7] = 8'h9d;
			8'h37 : d[0:7] = 8'h94;
			8'h38 : d[0:7] = 8'he3;
			8'h39 : d[0:7] = 8'hea;
			8'h3a : d[0:7] = 8'hf1;
			8'h3b : d[0:7] = 8'hf8;
			8'h3c : d[0:7] = 8'hc7;
			8'h3d : d[0:7] = 8'hce;
			8'h3e : d[0:7] = 8'hd5;
			8'h3f : d[0:7] = 8'hdc;
			8'h40 : d[0:7] = 8'h76;
			8'h41 : d[0:7] = 8'h7f;
			8'h42 : d[0:7] = 8'h64;
			8'h43 : d[0:7] = 8'h6d;
			8'h44 : d[0:7] = 8'h52;
			8'h45 : d[0:7] = 8'h5b;
			8'h46 : d[0:7] = 8'h40;
			8'h47 : d[0:7] = 8'h49;
			8'h48 : d[0:7] = 8'h3e;
			8'h49 : d[0:7] = 8'h37;
			8'h4a : d[0:7] = 8'h2c;
			8'h4b : d[0:7] = 8'h25;
			8'h4c : d[0:7] = 8'h1a;
			8'h4d : d[0:7] = 8'h13;
			8'h4e : d[0:7] = 8'h8;
			8'h4f : d[0:7] = 8'h1;
			8'h50 : d[0:7] = 8'he6;
			8'h51 : d[0:7] = 8'hef;
			8'h52 : d[0:7] = 8'hf4;
			8'h53 : d[0:7] = 8'hfd;
			8'h54 : d[0:7] = 8'hc2;
			8'h55 : d[0:7] = 8'hcb;
			8'h56 : d[0:7] = 8'hd0;
			8'h57 : d[0:7] = 8'hd9;
			8'h58 : d[0:7] = 8'hae;
			8'h59 : d[0:7] = 8'ha7;
			8'h5a : d[0:7] = 8'hbc;
			8'h5b : d[0:7] = 8'hb5;
			8'h5c : d[0:7] = 8'h8a;
			8'h5d : d[0:7] = 8'h83;
			8'h5e : d[0:7] = 8'h98;
			8'h5f : d[0:7] = 8'h91;
			8'h60 : d[0:7] = 8'h4d;
			8'h61 : d[0:7] = 8'h44;
			8'h62 : d[0:7] = 8'h5f;
			8'h63 : d[0:7] = 8'h56;
			8'h64 : d[0:7] = 8'h69;
			8'h65 : d[0:7] = 8'h60;
			8'h66 : d[0:7] = 8'h7b;
			8'h67 : d[0:7] = 8'h72;
			8'h68 : d[0:7] = 8'h5;
			8'h69 : d[0:7] = 8'hc;
			8'h6a : d[0:7] = 8'h17;
			8'h6b : d[0:7] = 8'h1e;
			8'h6c : d[0:7] = 8'h21;
			8'h6d : d[0:7] = 8'h28;
			8'h6e : d[0:7] = 8'h33;
			8'h6f : d[0:7] = 8'h3a;
			8'h70 : d[0:7] = 8'hdd;
			8'h71 : d[0:7] = 8'hd4;
			8'h72 : d[0:7] = 8'hcf;
			8'h73 : d[0:7] = 8'hc6;
			8'h74 : d[0:7] = 8'hf9;
			8'h75 : d[0:7] = 8'hf0;
			8'h76 : d[0:7] = 8'heb;
			8'h77 : d[0:7] = 8'he2;
			8'h78 : d[0:7] = 8'h95;
			8'h79 : d[0:7] = 8'h9c;
			8'h7a : d[0:7] = 8'h87;
			8'h7b : d[0:7] = 8'h8e;
			8'h7c : d[0:7] = 8'hb1;
			8'h7d : d[0:7] = 8'hb8;
			8'h7e : d[0:7] = 8'ha3;
			8'h7f : d[0:7] = 8'haa;
			8'h80 : d[0:7] = 8'hec;
			8'h81 : d[0:7] = 8'he5;
			8'h82 : d[0:7] = 8'hfe;
			8'h83 : d[0:7] = 8'hf7;
			8'h84 : d[0:7] = 8'hc8;
			8'h85 : d[0:7] = 8'hc1;
			8'h86 : d[0:7] = 8'hda;
			8'h87 : d[0:7] = 8'hd3;
			8'h88 : d[0:7] = 8'ha4;
			8'h89 : d[0:7] = 8'had;
			8'h8a : d[0:7] = 8'hb6;
			8'h8b : d[0:7] = 8'hbf;
			8'h8c : d[0:7] = 8'h80;
			8'h8d : d[0:7] = 8'h89;
			8'h8e : d[0:7] = 8'h92;
			8'h8f : d[0:7] = 8'h9b;
			8'h90 : d[0:7] = 8'h7c;
			8'h91 : d[0:7] = 8'h75;
			8'h92 : d[0:7] = 8'h6e;
			8'h93 : d[0:7] = 8'h67;
			8'h94 : d[0:7] = 8'h58;
			8'h95 : d[0:7] = 8'h51;
			8'h96 : d[0:7] = 8'h4a;
			8'h97 : d[0:7] = 8'h43;
			8'h98 : d[0:7] = 8'h34;
			8'h99 : d[0:7] = 8'h3d;
			8'h9a : d[0:7] = 8'h26;
			8'h9b : d[0:7] = 8'h2f;
			8'h9c : d[0:7] = 8'h10;
			8'h9d : d[0:7] = 8'h19;
			8'h9e : d[0:7] = 8'h2;
			8'h9f : d[0:7] = 8'hb;
			8'ha0 : d[0:7] = 8'hd7;
			8'ha1 : d[0:7] = 8'hde;
			8'ha2 : d[0:7] = 8'hc5;
			8'ha3 : d[0:7] = 8'hcc;
			8'ha4 : d[0:7] = 8'hf3;
			8'ha5 : d[0:7] = 8'hfa;
			8'ha6 : d[0:7] = 8'he1;
			8'ha7 : d[0:7] = 8'he8;
			8'ha8 : d[0:7] = 8'h9f;
			8'ha9 : d[0:7] = 8'h96;
			8'haa : d[0:7] = 8'h8d;
			8'hab : d[0:7] = 8'h84;
			8'hac : d[0:7] = 8'hbb;
			8'had : d[0:7] = 8'hb2;
			8'hae : d[0:7] = 8'ha9;
			8'haf : d[0:7] = 8'ha0;
			8'hb0 : d[0:7] = 8'h47;
			8'hb1 : d[0:7] = 8'h4e;
			8'hb2 : d[0:7] = 8'h55;
			8'hb3 : d[0:7] = 8'h5c;
			8'hb4 : d[0:7] = 8'h63;
			8'hb5 : d[0:7] = 8'h6a;
			8'hb6 : d[0:7] = 8'h71;
			8'hb7 : d[0:7] = 8'h78;
			8'hb8 : d[0:7] = 8'hf;
			8'hb9 : d[0:7] = 8'h6;
			8'hba : d[0:7] = 8'h1d;
			8'hbb : d[0:7] = 8'h14;
			8'hbc : d[0:7] = 8'h2b;
			8'hbd : d[0:7] = 8'h22;
			8'hbe : d[0:7] = 8'h39;
			8'hbf : d[0:7] = 8'h30;
			8'hc0 : d[0:7] = 8'h9a;
			8'hc1 : d[0:7] = 8'h93;
			8'hc2 : d[0:7] = 8'h88;
			8'hc3 : d[0:7] = 8'h81;
			8'hc4 : d[0:7] = 8'hbe;
			8'hc5 : d[0:7] = 8'hb7;
			8'hc6 : d[0:7] = 8'hac;
			8'hc7 : d[0:7] = 8'ha5;
			8'hc8 : d[0:7] = 8'hd2;
			8'hc9 : d[0:7] = 8'hdb;
			8'hca : d[0:7] = 8'hc0;
			8'hcb : d[0:7] = 8'hc9;
			8'hcc : d[0:7] = 8'hf6;
			8'hcd : d[0:7] = 8'hff;
			8'hce : d[0:7] = 8'he4;
			8'hcf : d[0:7] = 8'hed;
			8'hd0 : d[0:7] = 8'ha;
			8'hd1 : d[0:7] = 8'h3;
			8'hd2 : d[0:7] = 8'h18;
			8'hd3 : d[0:7] = 8'h11;
			8'hd4 : d[0:7] = 8'h2e;
			8'hd5 : d[0:7] = 8'h27;
			8'hd6 : d[0:7] = 8'h3c;
			8'hd7 : d[0:7] = 8'h35;
			8'hd8 : d[0:7] = 8'h42;
			8'hd9 : d[0:7] = 8'h4b;
			8'hda : d[0:7] = 8'h50;
			8'hdb : d[0:7] = 8'h59;
			8'hdc : d[0:7] = 8'h66;
			8'hdd : d[0:7] = 8'h6f;
			8'hde : d[0:7] = 8'h74;
			8'hdf : d[0:7] = 8'h7d;
			8'he0 : d[0:7] = 8'ha1;
			8'he1 : d[0:7] = 8'ha8;
			8'he2 : d[0:7] = 8'hb3;
			8'he3 : d[0:7] = 8'hba;
			8'he4 : d[0:7] = 8'h85;
			8'he5 : d[0:7] = 8'h8c;
			8'he6 : d[0:7] = 8'h97;
			8'he7 : d[0:7] = 8'h9e;
			8'he8 : d[0:7] = 8'he9;
			8'he9 : d[0:7] = 8'he0;
			8'hea : d[0:7] = 8'hfb;
			8'heb : d[0:7] = 8'hf2;
			8'hec : d[0:7] = 8'hcd;
			8'hed : d[0:7] = 8'hc4;
			8'hee : d[0:7] = 8'hdf;
			8'hef : d[0:7] = 8'hd6;
			8'hf0 : d[0:7] = 8'h31;
			8'hf1 : d[0:7] = 8'h38;
			8'hf2 : d[0:7] = 8'h23;
			8'hf3 : d[0:7] = 8'h2a;
			8'hf4 : d[0:7] = 8'h15;
			8'hf5 : d[0:7] = 8'h1c;
			8'hf6 : d[0:7] = 8'h7;
			8'hf7 : d[0:7] = 8'he;
			8'hf8 : d[0:7] = 8'h79;
			8'hf9 : d[0:7] = 8'h70;
			8'hfa : d[0:7] = 8'h6b;
			8'hfb : d[0:7] = 8'h62;
			8'hfc : d[0:7] = 8'h5d;
			8'hfd : d[0:7] = 8'h54;
			8'hfe : d[0:7] = 8'h4f;
			8'hff : d[0:7] = 8'h46;
        endcase
    end

    // Multiplication with 14
    always @(row[8:15]) begin
        case (row[8:15])
                        8'h0 : a[0:7] = 8'h0;
            8'h1 : a[0:7] = 8'he;
            8'h2 : a[0:7] = 8'h1c;
            8'h3 : a[0:7] = 8'h12;
            8'h4 : a[0:7] = 8'h38;
            8'h5 : a[0:7] = 8'h36;
            8'h6 : a[0:7] = 8'h24;
            8'h7 : a[0:7] = 8'h2a;
            8'h8 : a[0:7] = 8'h70;
            8'h9 : a[0:7] = 8'h7e;
            8'ha : a[0:7] = 8'h6c;
            8'hb : a[0:7] = 8'h62;
            8'hc : a[0:7] = 8'h48;
            8'hd : a[0:7] = 8'h46;
            8'he : a[0:7] = 8'h54;
            8'hf : a[0:7] = 8'h5a;
            8'h10 : a[0:7] = 8'he0;
            8'h11 : a[0:7] = 8'hee;
            8'h12 : a[0:7] = 8'hfc;
            8'h13 : a[0:7] = 8'hf2;
            8'h14 : a[0:7] = 8'hd8;
            8'h15 : a[0:7] = 8'hd6;
            8'h16 : a[0:7] = 8'hc4;
            8'h17 : a[0:7] = 8'hca;
            8'h18 : a[0:7] = 8'h90;
            8'h19 : a[0:7] = 8'h9e;
            8'h1a : a[0:7] = 8'h8c;
            8'h1b : a[0:7] = 8'h82;
            8'h1c : a[0:7] = 8'ha8;
            8'h1d : a[0:7] = 8'ha6;
            8'h1e : a[0:7] = 8'hb4;
            8'h1f : a[0:7] = 8'hba;
            8'h20 : a[0:7] = 8'hdb;
            8'h21 : a[0:7] = 8'hd5;
            8'h22 : a[0:7] = 8'hc7;
            8'h23 : a[0:7] = 8'hc9;
            8'h24 : a[0:7] = 8'he3;
            8'h25 : a[0:7] = 8'hed;
            8'h26 : a[0:7] = 8'hff;
            8'h27 : a[0:7] = 8'hf1;
            8'h28 : a[0:7] = 8'hab;
            8'h29 : a[0:7] = 8'ha5;
            8'h2a : a[0:7] = 8'hb7;
            8'h2b : a[0:7] = 8'hb9;
            8'h2c : a[0:7] = 8'h93;
            8'h2d : a[0:7] = 8'h9d;
            8'h2e : a[0:7] = 8'h8f;
            8'h2f : a[0:7] = 8'h81;
            8'h30 : a[0:7] = 8'h3b;
            8'h31 : a[0:7] = 8'h35;
            8'h32 : a[0:7] = 8'h27;
            8'h33 : a[0:7] = 8'h29;
            8'h34 : a[0:7] = 8'h3;
            8'h35 : a[0:7] = 8'hd;
            8'h36 : a[0:7] = 8'h1f;
            8'h37 : a[0:7] = 8'h11;
            8'h38 : a[0:7] = 8'h4b;
            8'h39 : a[0:7] = 8'h45;
            8'h3a : a[0:7] = 8'h57;
            8'h3b : a[0:7] = 8'h59;
            8'h3c : a[0:7] = 8'h73;
            8'h3d : a[0:7] = 8'h7d;
            8'h3e : a[0:7] = 8'h6f;
            8'h3f : a[0:7] = 8'h61;
            8'h40 : a[0:7] = 8'had;
            8'h41 : a[0:7] = 8'ha3;
            8'h42 : a[0:7] = 8'hb1;
            8'h43 : a[0:7] = 8'hbf;
            8'h44 : a[0:7] = 8'h95;
            8'h45 : a[0:7] = 8'h9b;
            8'h46 : a[0:7] = 8'h89;
            8'h47 : a[0:7] = 8'h87;
            8'h48 : a[0:7] = 8'hdd;
            8'h49 : a[0:7] = 8'hd3;
            8'h4a : a[0:7] = 8'hc1;
            8'h4b : a[0:7] = 8'hcf;
            8'h4c : a[0:7] = 8'he5;
            8'h4d : a[0:7] = 8'heb;
            8'h4e : a[0:7] = 8'hf9;
            8'h4f : a[0:7] = 8'hf7;
            8'h50 : a[0:7] = 8'h4d;
            8'h51 : a[0:7] = 8'h43;
            8'h52 : a[0:7] = 8'h51;
            8'h53 : a[0:7] = 8'h5f;
            8'h54 : a[0:7] = 8'h75;
            8'h55 : a[0:7] = 8'h7b;
            8'h56 : a[0:7] = 8'h69;
            8'h57 : a[0:7] = 8'h67;
            8'h58 : a[0:7] = 8'h3d;
            8'h59 : a[0:7] = 8'h33;
            8'h5a : a[0:7] = 8'h21;
            8'h5b : a[0:7] = 8'h2f;
            8'h5c : a[0:7] = 8'h5;
            8'h5d : a[0:7] = 8'hb;
            8'h5e : a[0:7] = 8'h19;
            8'h5f : a[0:7] = 8'h17;
            8'h60 : a[0:7] = 8'h76;
            8'h61 : a[0:7] = 8'h78;
            8'h62 : a[0:7] = 8'h6a;
            8'h63 : a[0:7] = 8'h64;
            8'h64 : a[0:7] = 8'h4e;
            8'h65 : a[0:7] = 8'h40;
            8'h66 : a[0:7] = 8'h52;
            8'h67 : a[0:7] = 8'h5c;
            8'h68 : a[0:7] = 8'h6;
            8'h69 : a[0:7] = 8'h8;
            8'h6a : a[0:7] = 8'h1a;
            8'h6b : a[0:7] = 8'h14;
            8'h6c : a[0:7] = 8'h3e;
            8'h6d : a[0:7] = 8'h30;
            8'h6e : a[0:7] = 8'h22;
            8'h6f : a[0:7] = 8'h2c;
            8'h70 : a[0:7] = 8'h96;
            8'h71 : a[0:7] = 8'h98;
            8'h72 : a[0:7] = 8'h8a;
            8'h73 : a[0:7] = 8'h84;
            8'h74 : a[0:7] = 8'hae;
            8'h75 : a[0:7] = 8'ha0;
            8'h76 : a[0:7] = 8'hb2;
            8'h77 : a[0:7] = 8'hbc;
            8'h78 : a[0:7] = 8'he6;
            8'h79 : a[0:7] = 8'he8;
            8'h7a : a[0:7] = 8'hfa;
            8'h7b : a[0:7] = 8'hf4;
            8'h7c : a[0:7] = 8'hde;
            8'h7d : a[0:7] = 8'hd0;
            8'h7e : a[0:7] = 8'hc2;
            8'h7f : a[0:7] = 8'hcc;
            8'h80 : a[0:7] = 8'h41;
            8'h81 : a[0:7] = 8'h4f;
            8'h82 : a[0:7] = 8'h5d;
            8'h83 : a[0:7] = 8'h53;
            8'h84 : a[0:7] = 8'h79;
            8'h85 : a[0:7] = 8'h77;
            8'h86 : a[0:7] = 8'h65;
            8'h87 : a[0:7] = 8'h6b;
            8'h88 : a[0:7] = 8'h31;
            8'h89 : a[0:7] = 8'h3f;
            8'h8a : a[0:7] = 8'h2d;
            8'h8b : a[0:7] = 8'h23;
            8'h8c : a[0:7] = 8'h9;
            8'h8d : a[0:7] = 8'h7;
            8'h8e : a[0:7] = 8'h15;
            8'h8f : a[0:7] = 8'h1b;
            8'h90 : a[0:7] = 8'ha1;
            8'h91 : a[0:7] = 8'haf;
            8'h92 : a[0:7] = 8'hbd;
            8'h93 : a[0:7] = 8'hb3;
            8'h94 : a[0:7] = 8'h99;
            8'h95 : a[0:7] = 8'h97;
            8'h96 : a[0:7] = 8'h85;
            8'h97 : a[0:7] = 8'h8b;
            8'h98 : a[0:7] = 8'hd1;
            8'h99 : a[0:7] = 8'hdf;
            8'h9a : a[0:7] = 8'hcd;
            8'h9b : a[0:7] = 8'hc3;
            8'h9c : a[0:7] = 8'he9;
            8'h9d : a[0:7] = 8'he7;
            8'h9e : a[0:7] = 8'hf5;
            8'h9f : a[0:7] = 8'hfb;
            8'ha0 : a[0:7] = 8'h9a;
            8'ha1 : a[0:7] = 8'h94;
            8'ha2 : a[0:7] = 8'h86;
            8'ha3 : a[0:7] = 8'h88;
            8'ha4 : a[0:7] = 8'ha2;
            8'ha5 : a[0:7] = 8'hac;
            8'ha6 : a[0:7] = 8'hbe;
            8'ha7 : a[0:7] = 8'hb0;
            8'ha8 : a[0:7] = 8'hea;
            8'ha9 : a[0:7] = 8'he4;
            8'haa : a[0:7] = 8'hf6;
            8'hab : a[0:7] = 8'hf8;
            8'hac : a[0:7] = 8'hd2;
            8'had : a[0:7] = 8'hdc;
            8'hae : a[0:7] = 8'hce;
            8'haf : a[0:7] = 8'hc0;
            8'hb0 : a[0:7] = 8'h7a;
            8'hb1 : a[0:7] = 8'h74;
            8'hb2 : a[0:7] = 8'h66;
            8'hb3 : a[0:7] = 8'h68;
            8'hb4 : a[0:7] = 8'h42;
            8'hb5 : a[0:7] = 8'h4c;
            8'hb6 : a[0:7] = 8'h5e;
            8'hb7 : a[0:7] = 8'h50;
            8'hb8 : a[0:7] = 8'ha;
            8'hb9 : a[0:7] = 8'h4;
            8'hba : a[0:7] = 8'h16;
            8'hbb : a[0:7] = 8'h18;
            8'hbc : a[0:7] = 8'h32;
            8'hbd : a[0:7] = 8'h3c;
            8'hbe : a[0:7] = 8'h2e;
            8'hbf : a[0:7] = 8'h20;
            8'hc0 : a[0:7] = 8'hec;
            8'hc1 : a[0:7] = 8'he2;
            8'hc2 : a[0:7] = 8'hf0;
            8'hc3 : a[0:7] = 8'hfe;
            8'hc4 : a[0:7] = 8'hd4;
            8'hc5 : a[0:7] = 8'hda;
            8'hc6 : a[0:7] = 8'hc8;
            8'hc7 : a[0:7] = 8'hc6;
            8'hc8 : a[0:7] = 8'h9c;
            8'hc9 : a[0:7] = 8'h92;
            8'hca : a[0:7] = 8'h80;
            8'hcb : a[0:7] = 8'h8e;
            8'hcc : a[0:7] = 8'ha4;
            8'hcd : a[0:7] = 8'haa;
            8'hce : a[0:7] = 8'hb8;
            8'hcf : a[0:7] = 8'hb6;
            8'hd0 : a[0:7] = 8'hc;
            8'hd1 : a[0:7] = 8'h2;
            8'hd2 : a[0:7] = 8'h10;
            8'hd3 : a[0:7] = 8'h1e;
            8'hd4 : a[0:7] = 8'h34;
            8'hd5 : a[0:7] = 8'h3a;
            8'hd6 : a[0:7] = 8'h28;
            8'hd7 : a[0:7] = 8'h26;
            8'hd8 : a[0:7] = 8'h7c;
            8'hd9 : a[0:7] = 8'h72;
            8'hda : a[0:7] = 8'h60;
            8'hdb : a[0:7] = 8'h6e;
            8'hdc : a[0:7] = 8'h44;
            8'hdd : a[0:7] = 8'h4a;
            8'hde : a[0:7] = 8'h58;
            8'hdf : a[0:7] = 8'h56;
            8'he0 : a[0:7] = 8'h37;
            8'he1 : a[0:7] = 8'h39;
            8'he2 : a[0:7] = 8'h2b;
            8'he3 : a[0:7] = 8'h25;
            8'he4 : a[0:7] = 8'hf;
            8'he5 : a[0:7] = 8'h1;
            8'he6 : a[0:7] = 8'h13;
            8'he7 : a[0:7] = 8'h1d;
            8'he8 : a[0:7] = 8'h47;
            8'he9 : a[0:7] = 8'h49;
            8'hea : a[0:7] = 8'h5b;
            8'heb : a[0:7] = 8'h55;
            8'hec : a[0:7] = 8'h7f;
            8'hed : a[0:7] = 8'h71;
            8'hee : a[0:7] = 8'h63;
            8'hef : a[0:7] = 8'h6d;
            8'hf0 : a[0:7] = 8'hd7;
            8'hf1 : a[0:7] = 8'hd9;
            8'hf2 : a[0:7] = 8'hcb;
            8'hf3 : a[0:7] = 8'hc5;
            8'hf4 : a[0:7] = 8'hef;
            8'hf5 : a[0:7] = 8'he1;
            8'hf6 : a[0:7] = 8'hf3;
            8'hf7 : a[0:7] = 8'hfd;
            8'hf8 : a[0:7] = 8'ha7;
            8'hf9 : a[0:7] = 8'ha9;
            8'hfa : a[0:7] = 8'hbb;
            8'hfb : a[0:7] = 8'hb5;
            8'hfc : a[0:7] = 8'h9f;
            8'hfd : a[0:7] = 8'h91;
            8'hfe : a[0:7] = 8'h83;
            8'hff : a[0:7] = 8'h8d;
        endcase
    end

    // Multiplication with 11
    always @(row[16:23]) begin
        case (row[16:23])
			            8'h0 : b[0:7] = 8'h0;
            8'h1 : b[0:7] = 8'hb;
            8'h2 : b[0:7] = 8'h16;
            8'h3 : b[0:7] = 8'h1d;
            8'h4 : b[0:7] = 8'h2c;
            8'h5 : b[0:7] = 8'h27;
            8'h6 : b[0:7] = 8'h3a;
            8'h7 : b[0:7] = 8'h31;
            8'h8 : b[0:7] = 8'h58;
            8'h9 : b[0:7] = 8'h53;
            8'ha : b[0:7] = 8'h4e;
            8'hb : b[0:7] = 8'h45;
            8'hc : b[0:7] = 8'h74;
            8'hd : b[0:7] = 8'h7f;
            8'he : b[0:7] = 8'h62;
            8'hf : b[0:7] = 8'h69;
            8'h10 : b[0:7] = 8'hb0;
            8'h11 : b[0:7] = 8'hbb;
            8'h12 : b[0:7] = 8'ha6;
            8'h13 : b[0:7] = 8'had;
            8'h14 : b[0:7] = 8'h9c;
            8'h15 : b[0:7] = 8'h97;
            8'h16 : b[0:7] = 8'h8a;
            8'h17 : b[0:7] = 8'h81;
            8'h18 : b[0:7] = 8'he8;
            8'h19 : b[0:7] = 8'he3;
            8'h1a : b[0:7] = 8'hfe;
            8'h1b : b[0:7] = 8'hf5;
            8'h1c : b[0:7] = 8'hc4;
            8'h1d : b[0:7] = 8'hcf;
            8'h1e : b[0:7] = 8'hd2;
            8'h1f : b[0:7] = 8'hd9;
            8'h20 : b[0:7] = 8'h7b;
            8'h21 : b[0:7] = 8'h70;
            8'h22 : b[0:7] = 8'h6d;
            8'h23 : b[0:7] = 8'h66;
            8'h24 : b[0:7] = 8'h57;
            8'h25 : b[0:7] = 8'h5c;
            8'h26 : b[0:7] = 8'h41;
            8'h27 : b[0:7] = 8'h4a;
            8'h28 : b[0:7] = 8'h23;
            8'h29 : b[0:7] = 8'h28;
            8'h2a : b[0:7] = 8'h35;
            8'h2b : b[0:7] = 8'h3e;
            8'h2c : b[0:7] = 8'hf;
            8'h2d : b[0:7] = 8'h4;
            8'h2e : b[0:7] = 8'h19;
            8'h2f : b[0:7] = 8'h12;
            8'h30 : b[0:7] = 8'hcb;
            8'h31 : b[0:7] = 8'hc0;
            8'h32 : b[0:7] = 8'hdd;
            8'h33 : b[0:7] = 8'hd6;
            8'h34 : b[0:7] = 8'he7;
            8'h35 : b[0:7] = 8'hec;
            8'h36 : b[0:7] = 8'hf1;
            8'h37 : b[0:7] = 8'hfa;
            8'h38 : b[0:7] = 8'h93;
            8'h39 : b[0:7] = 8'h98;
            8'h3a : b[0:7] = 8'h85;
            8'h3b : b[0:7] = 8'h8e;
            8'h3c : b[0:7] = 8'hbf;
            8'h3d : b[0:7] = 8'hb4;
            8'h3e : b[0:7] = 8'ha9;
            8'h3f : b[0:7] = 8'ha2;
            8'h40 : b[0:7] = 8'hf6;
            8'h41 : b[0:7] = 8'hfd;
            8'h42 : b[0:7] = 8'he0;
            8'h43 : b[0:7] = 8'heb;
            8'h44 : b[0:7] = 8'hda;
            8'h45 : b[0:7] = 8'hd1;
            8'h46 : b[0:7] = 8'hcc;
            8'h47 : b[0:7] = 8'hc7;
            8'h48 : b[0:7] = 8'hae;
            8'h49 : b[0:7] = 8'ha5;
            8'h4a : b[0:7] = 8'hb8;
            8'h4b : b[0:7] = 8'hb3;
            8'h4c : b[0:7] = 8'h82;
            8'h4d : b[0:7] = 8'h89;
            8'h4e : b[0:7] = 8'h94;
            8'h4f : b[0:7] = 8'h9f;
            8'h50 : b[0:7] = 8'h46;
            8'h51 : b[0:7] = 8'h4d;
            8'h52 : b[0:7] = 8'h50;
            8'h53 : b[0:7] = 8'h5b;
            8'h54 : b[0:7] = 8'h6a;
            8'h55 : b[0:7] = 8'h61;
            8'h56 : b[0:7] = 8'h7c;
            8'h57 : b[0:7] = 8'h77;
            8'h58 : b[0:7] = 8'h1e;
            8'h59 : b[0:7] = 8'h15;
            8'h5a : b[0:7] = 8'h8;
            8'h5b : b[0:7] = 8'h3;
            8'h5c : b[0:7] = 8'h32;
            8'h5d : b[0:7] = 8'h39;
            8'h5e : b[0:7] = 8'h24;
            8'h5f : b[0:7] = 8'h2f;
            8'h60 : b[0:7] = 8'h8d;
            8'h61 : b[0:7] = 8'h86;
            8'h62 : b[0:7] = 8'h9b;
            8'h63 : b[0:7] = 8'h90;
            8'h64 : b[0:7] = 8'ha1;
            8'h65 : b[0:7] = 8'haa;
            8'h66 : b[0:7] = 8'hb7;
            8'h67 : b[0:7] = 8'hbc;
            8'h68 : b[0:7] = 8'hd5;
            8'h69 : b[0:7] = 8'hde;
            8'h6a : b[0:7] = 8'hc3;
            8'h6b : b[0:7] = 8'hc8;
            8'h6c : b[0:7] = 8'hf9;
            8'h6d : b[0:7] = 8'hf2;
            8'h6e : b[0:7] = 8'hef;
            8'h6f : b[0:7] = 8'he4;
            8'h70 : b[0:7] = 8'h3d;
            8'h71 : b[0:7] = 8'h36;
            8'h72 : b[0:7] = 8'h2b;
            8'h73 : b[0:7] = 8'h20;
            8'h74 : b[0:7] = 8'h11;
            8'h75 : b[0:7] = 8'h1a;
            8'h76 : b[0:7] = 8'h7;
            8'h77 : b[0:7] = 8'hc;
            8'h78 : b[0:7] = 8'h65;
            8'h79 : b[0:7] = 8'h6e;
            8'h7a : b[0:7] = 8'h73;
            8'h7b : b[0:7] = 8'h78;
            8'h7c : b[0:7] = 8'h49;
            8'h7d : b[0:7] = 8'h42;
            8'h7e : b[0:7] = 8'h5f;
            8'h7f : b[0:7] = 8'h54;
            8'h80 : b[0:7] = 8'hf7;
            8'h81 : b[0:7] = 8'hfc;
            8'h82 : b[0:7] = 8'he1;
            8'h83 : b[0:7] = 8'hea;
            8'h84 : b[0:7] = 8'hdb;
            8'h85 : b[0:7] = 8'hd0;
            8'h86 : b[0:7] = 8'hcd;
            8'h87 : b[0:7] = 8'hc6;
            8'h88 : b[0:7] = 8'haf;
            8'h89 : b[0:7] = 8'ha4;
            8'h8a : b[0:7] = 8'hb9;
            8'h8b : b[0:7] = 8'hb2;
            8'h8c : b[0:7] = 8'h83;
            8'h8d : b[0:7] = 8'h88;
            8'h8e : b[0:7] = 8'h95;
            8'h8f : b[0:7] = 8'h9e;
            8'h90 : b[0:7] = 8'h47;
            8'h91 : b[0:7] = 8'h4c;
            8'h92 : b[0:7] = 8'h51;
            8'h93 : b[0:7] = 8'h5a;
            8'h94 : b[0:7] = 8'h6b;
            8'h95 : b[0:7] = 8'h60;
            8'h96 : b[0:7] = 8'h7d;
            8'h97 : b[0:7] = 8'h76;
            8'h98 : b[0:7] = 8'h1f;
            8'h99 : b[0:7] = 8'h14;
            8'h9a : b[0:7] = 8'h9;
            8'h9b : b[0:7] = 8'h2;
            8'h9c : b[0:7] = 8'h33;
            8'h9d : b[0:7] = 8'h38;
            8'h9e : b[0:7] = 8'h25;
            8'h9f : b[0:7] = 8'h2e;
            8'ha0 : b[0:7] = 8'h8c;
            8'ha1 : b[0:7] = 8'h87;
            8'ha2 : b[0:7] = 8'h9a;
            8'ha3 : b[0:7] = 8'h91;
            8'ha4 : b[0:7] = 8'ha0;
            8'ha5 : b[0:7] = 8'hab;
            8'ha6 : b[0:7] = 8'hb6;
            8'ha7 : b[0:7] = 8'hbd;
            8'ha8 : b[0:7] = 8'hd4;
            8'ha9 : b[0:7] = 8'hdf;
            8'haa : b[0:7] = 8'hc2;
            8'hab : b[0:7] = 8'hc9;
            8'hac : b[0:7] = 8'hf8;
            8'had : b[0:7] = 8'hf3;
            8'hae : b[0:7] = 8'hee;
            8'haf : b[0:7] = 8'he5;
            8'hb0 : b[0:7] = 8'h3c;
            8'hb1 : b[0:7] = 8'h37;
            8'hb2 : b[0:7] = 8'h2a;
            8'hb3 : b[0:7] = 8'h21;
            8'hb4 : b[0:7] = 8'h10;
            8'hb5 : b[0:7] = 8'h1b;
            8'hb6 : b[0:7] = 8'h6;
            8'hb7 : b[0:7] = 8'hd;
            8'hb8 : b[0:7] = 8'h64;
            8'hb9 : b[0:7] = 8'h6f;
            8'hba : b[0:7] = 8'h72;
            8'hbb : b[0:7] = 8'h79;
            8'hbc : b[0:7] = 8'h48;
            8'hbd : b[0:7] = 8'h43;
            8'hbe : b[0:7] = 8'h5e;
            8'hbf : b[0:7] = 8'h55;
            8'hc0 : b[0:7] = 8'h1;
            8'hc1 : b[0:7] = 8'ha;
            8'hc2 : b[0:7] = 8'h17;
            8'hc3 : b[0:7] = 8'h1c;
            8'hc4 : b[0:7] = 8'h2d;
            8'hc5 : b[0:7] = 8'h26;
            8'hc6 : b[0:7] = 8'h3b;
            8'hc7 : b[0:7] = 8'h30;
            8'hc8 : b[0:7] = 8'h59;
            8'hc9 : b[0:7] = 8'h52;
            8'hca : b[0:7] = 8'h4f;
            8'hcb : b[0:7] = 8'h44;
            8'hcc : b[0:7] = 8'h75;
            8'hcd : b[0:7] = 8'h7e;
            8'hce : b[0:7] = 8'h63;
            8'hcf : b[0:7] = 8'h68;
            8'hd0 : b[0:7] = 8'hb1;
            8'hd1 : b[0:7] = 8'hba;
            8'hd2 : b[0:7] = 8'ha7;
            8'hd3 : b[0:7] = 8'hac;
            8'hd4 : b[0:7] = 8'h9d;
            8'hd5 : b[0:7] = 8'h96;
            8'hd6 : b[0:7] = 8'h8b;
            8'hd7 : b[0:7] = 8'h80;
            8'hd8 : b[0:7] = 8'he9;
            8'hd9 : b[0:7] = 8'he2;
            8'hda : b[0:7] = 8'hff;
            8'hdb : b[0:7] = 8'hf4;
            8'hdc : b[0:7] = 8'hc5;
            8'hdd : b[0:7] = 8'hce;
            8'hde : b[0:7] = 8'hd3;
            8'hdf : b[0:7] = 8'hd8;
            8'he0 : b[0:7] = 8'h7a;
            8'he1 : b[0:7] = 8'h71;
            8'he2 : b[0:7] = 8'h6c;
            8'he3 : b[0:7] = 8'h67;
            8'he4 : b[0:7] = 8'h56;
            8'he5 : b[0:7] = 8'h5d;
            8'he6 : b[0:7] = 8'h40;
            8'he7 : b[0:7] = 8'h4b;
            8'he8 : b[0:7] = 8'h22;
            8'he9 : b[0:7] = 8'h29;
            8'hea : b[0:7] = 8'h34;
            8'heb : b[0:7] = 8'h3f;
            8'hec : b[0:7] = 8'he;
            8'hed : b[0:7] = 8'h5;
            8'hee : b[0:7] = 8'h18;
            8'hef : b[0:7] = 8'h13;
            8'hf0 : b[0:7] = 8'hca;
            8'hf1 : b[0:7] = 8'hc1;
            8'hf2 : b[0:7] = 8'hdc;
            8'hf3 : b[0:7] = 8'hd7;
            8'hf4 : b[0:7] = 8'he6;
            8'hf5 : b[0:7] = 8'hed;
            8'hf6 : b[0:7] = 8'hf0;
            8'hf7 : b[0:7] = 8'hfb;
            8'hf8 : b[0:7] = 8'h92;
            8'hf9 : b[0:7] = 8'h99;
            8'hfa : b[0:7] = 8'h84;
            8'hfb : b[0:7] = 8'h8f;
            8'hfc : b[0:7] = 8'hbe;
            8'hfd : b[0:7] = 8'hb5;
            8'hfe : b[0:7] = 8'ha8;
            8'hff : b[0:7] = 8'ha3;
        endcase
    end

    // Multiplication with 13
    always @(row[24:31]) begin
        case (row[24:31])
						8'h0 : c[0:7] = 8'h0;
			8'h1 : c[0:7] = 8'hd;
			8'h2 : c[0:7] = 8'h1a;
			8'h3 : c[0:7] = 8'h17;
			8'h4 : c[0:7] = 8'h34;
			8'h5 : c[0:7] = 8'h39;
			8'h6 : c[0:7] = 8'h2e;
			8'h7 : c[0:7] = 8'h23;
			8'h8 : c[0:7] = 8'h68;
			8'h9 : c[0:7] = 8'h65;
			8'ha : c[0:7] = 8'h72;
			8'hb : c[0:7] = 8'h7f;
			8'hc : c[0:7] = 8'h5c;
			8'hd : c[0:7] = 8'h51;
			8'he : c[0:7] = 8'h46;
			8'hf : c[0:7] = 8'h4b;
			8'h10 : c[0:7] = 8'hd0;
			8'h11 : c[0:7] = 8'hdd;
			8'h12 : c[0:7] = 8'hca;
			8'h13 : c[0:7] = 8'hc7;
			8'h14 : c[0:7] = 8'he4;
			8'h15 : c[0:7] = 8'he9;
			8'h16 : c[0:7] = 8'hfe;
			8'h17 : c[0:7] = 8'hf3;
			8'h18 : c[0:7] = 8'hb8;
			8'h19 : c[0:7] = 8'hb5;
			8'h1a : c[0:7] = 8'ha2;
			8'h1b : c[0:7] = 8'haf;
			8'h1c : c[0:7] = 8'h8c;
			8'h1d : c[0:7] = 8'h81;
			8'h1e : c[0:7] = 8'h96;
			8'h1f : c[0:7] = 8'h9b;
			8'h20 : c[0:7] = 8'hbb;
			8'h21 : c[0:7] = 8'hb6;
			8'h22 : c[0:7] = 8'ha1;
			8'h23 : c[0:7] = 8'hac;
			8'h24 : c[0:7] = 8'h8f;
			8'h25 : c[0:7] = 8'h82;
			8'h26 : c[0:7] = 8'h95;
			8'h27 : c[0:7] = 8'h98;
			8'h28 : c[0:7] = 8'hd3;
			8'h29 : c[0:7] = 8'hde;
			8'h2a : c[0:7] = 8'hc9;
			8'h2b : c[0:7] = 8'hc4;
			8'h2c : c[0:7] = 8'he7;
			8'h2d : c[0:7] = 8'hea;
			8'h2e : c[0:7] = 8'hfd;
			8'h2f : c[0:7] = 8'hf0;
			8'h30 : c[0:7] = 8'h6b;
			8'h31 : c[0:7] = 8'h66;
			8'h32 : c[0:7] = 8'h71;
			8'h33 : c[0:7] = 8'h7c;
			8'h34 : c[0:7] = 8'h5f;
			8'h35 : c[0:7] = 8'h52;
			8'h36 : c[0:7] = 8'h45;
			8'h37 : c[0:7] = 8'h48;
			8'h38 : c[0:7] = 8'h3;
			8'h39 : c[0:7] = 8'he;
			8'h3a : c[0:7] = 8'h19;
			8'h3b : c[0:7] = 8'h14;
			8'h3c : c[0:7] = 8'h37;
			8'h3d : c[0:7] = 8'h3a;
			8'h3e : c[0:7] = 8'h2d;
			8'h3f : c[0:7] = 8'h20;
			8'h40 : c[0:7] = 8'h6d;
			8'h41 : c[0:7] = 8'h60;
			8'h42 : c[0:7] = 8'h77;
			8'h43 : c[0:7] = 8'h7a;
			8'h44 : c[0:7] = 8'h59;
			8'h45 : c[0:7] = 8'h54;
			8'h46 : c[0:7] = 8'h43;
			8'h47 : c[0:7] = 8'h4e;
			8'h48 : c[0:7] = 8'h5;
			8'h49 : c[0:7] = 8'h8;
			8'h4a : c[0:7] = 8'h1f;
			8'h4b : c[0:7] = 8'h12;
			8'h4c : c[0:7] = 8'h31;
			8'h4d : c[0:7] = 8'h3c;
			8'h4e : c[0:7] = 8'h2b;
			8'h4f : c[0:7] = 8'h26;
			8'h50 : c[0:7] = 8'hbd;
			8'h51 : c[0:7] = 8'hb0;
			8'h52 : c[0:7] = 8'ha7;
			8'h53 : c[0:7] = 8'haa;
			8'h54 : c[0:7] = 8'h89;
			8'h55 : c[0:7] = 8'h84;
			8'h56 : c[0:7] = 8'h93;
			8'h57 : c[0:7] = 8'h9e;
			8'h58 : c[0:7] = 8'hd5;
			8'h59 : c[0:7] = 8'hd8;
			8'h5a : c[0:7] = 8'hcf;
			8'h5b : c[0:7] = 8'hc2;
			8'h5c : c[0:7] = 8'he1;
			8'h5d : c[0:7] = 8'hec;
			8'h5e : c[0:7] = 8'hfb;
			8'h5f : c[0:7] = 8'hf6;
			8'h60 : c[0:7] = 8'hd6;
			8'h61 : c[0:7] = 8'hdb;
			8'h62 : c[0:7] = 8'hcc;
			8'h63 : c[0:7] = 8'hc1;
			8'h64 : c[0:7] = 8'he2;
			8'h65 : c[0:7] = 8'hef;
			8'h66 : c[0:7] = 8'hf8;
			8'h67 : c[0:7] = 8'hf5;
			8'h68 : c[0:7] = 8'hbe;
			8'h69 : c[0:7] = 8'hb3;
			8'h6a : c[0:7] = 8'ha4;
			8'h6b : c[0:7] = 8'ha9;
			8'h6c : c[0:7] = 8'h8a;
			8'h6d : c[0:7] = 8'h87;
			8'h6e : c[0:7] = 8'h90;
			8'h6f : c[0:7] = 8'h9d;
			8'h70 : c[0:7] = 8'h6;
			8'h71 : c[0:7] = 8'hb;
			8'h72 : c[0:7] = 8'h1c;
			8'h73 : c[0:7] = 8'h11;
			8'h74 : c[0:7] = 8'h32;
			8'h75 : c[0:7] = 8'h3f;
			8'h76 : c[0:7] = 8'h28;
			8'h77 : c[0:7] = 8'h25;
			8'h78 : c[0:7] = 8'h6e;
			8'h79 : c[0:7] = 8'h63;
			8'h7a : c[0:7] = 8'h74;
			8'h7b : c[0:7] = 8'h79;
			8'h7c : c[0:7] = 8'h5a;
			8'h7d : c[0:7] = 8'h57;
			8'h7e : c[0:7] = 8'h40;
			8'h7f : c[0:7] = 8'h4d;
			8'h80 : c[0:7] = 8'hda;
			8'h81 : c[0:7] = 8'hd7;
			8'h82 : c[0:7] = 8'hc0;
			8'h83 : c[0:7] = 8'hcd;
			8'h84 : c[0:7] = 8'hee;
			8'h85 : c[0:7] = 8'he3;
			8'h86 : c[0:7] = 8'hf4;
			8'h87 : c[0:7] = 8'hf9;
			8'h88 : c[0:7] = 8'hb2;
			8'h89 : c[0:7] = 8'hbf;
			8'h8a : c[0:7] = 8'ha8;
			8'h8b : c[0:7] = 8'ha5;
			8'h8c : c[0:7] = 8'h86;
			8'h8d : c[0:7] = 8'h8b;
			8'h8e : c[0:7] = 8'h9c;
			8'h8f : c[0:7] = 8'h91;
			8'h90 : c[0:7] = 8'ha;
			8'h91 : c[0:7] = 8'h7;
			8'h92 : c[0:7] = 8'h10;
			8'h93 : c[0:7] = 8'h1d;
			8'h94 : c[0:7] = 8'h3e;
			8'h95 : c[0:7] = 8'h33;
			8'h96 : c[0:7] = 8'h24;
			8'h97 : c[0:7] = 8'h29;
			8'h98 : c[0:7] = 8'h62;
			8'h99 : c[0:7] = 8'h6f;
			8'h9a : c[0:7] = 8'h78;
			8'h9b : c[0:7] = 8'h75;
			8'h9c : c[0:7] = 8'h56;
			8'h9d : c[0:7] = 8'h5b;
			8'h9e : c[0:7] = 8'h4c;
			8'h9f : c[0:7] = 8'h41;
			8'ha0 : c[0:7] = 8'h61;
			8'ha1 : c[0:7] = 8'h6c;
			8'ha2 : c[0:7] = 8'h7b;
			8'ha3 : c[0:7] = 8'h76;
			8'ha4 : c[0:7] = 8'h55;
			8'ha5 : c[0:7] = 8'h58;
			8'ha6 : c[0:7] = 8'h4f;
			8'ha7 : c[0:7] = 8'h42;
			8'ha8 : c[0:7] = 8'h9;
			8'ha9 : c[0:7] = 8'h4;
			8'haa : c[0:7] = 8'h13;
			8'hab : c[0:7] = 8'h1e;
			8'hac : c[0:7] = 8'h3d;
			8'had : c[0:7] = 8'h30;
			8'hae : c[0:7] = 8'h27;
			8'haf : c[0:7] = 8'h2a;
			8'hb0 : c[0:7] = 8'hb1;
			8'hb1 : c[0:7] = 8'hbc;
			8'hb2 : c[0:7] = 8'hab;
			8'hb3 : c[0:7] = 8'ha6;
			8'hb4 : c[0:7] = 8'h85;
			8'hb5 : c[0:7] = 8'h88;
			8'hb6 : c[0:7] = 8'h9f;
			8'hb7 : c[0:7] = 8'h92;
			8'hb8 : c[0:7] = 8'hd9;
			8'hb9 : c[0:7] = 8'hd4;
			8'hba : c[0:7] = 8'hc3;
			8'hbb : c[0:7] = 8'hce;
			8'hbc : c[0:7] = 8'hed;
			8'hbd : c[0:7] = 8'he0;
			8'hbe : c[0:7] = 8'hf7;
			8'hbf : c[0:7] = 8'hfa;
			8'hc0 : c[0:7] = 8'hb7;
			8'hc1 : c[0:7] = 8'hba;
			8'hc2 : c[0:7] = 8'had;
			8'hc3 : c[0:7] = 8'ha0;
			8'hc4 : c[0:7] = 8'h83;
			8'hc5 : c[0:7] = 8'h8e;
			8'hc6 : c[0:7] = 8'h99;
			8'hc7 : c[0:7] = 8'h94;
			8'hc8 : c[0:7] = 8'hdf;
			8'hc9 : c[0:7] = 8'hd2;
			8'hca : c[0:7] = 8'hc5;
			8'hcb : c[0:7] = 8'hc8;
			8'hcc : c[0:7] = 8'heb;
			8'hcd : c[0:7] = 8'he6;
			8'hce : c[0:7] = 8'hf1;
			8'hcf : c[0:7] = 8'hfc;
			8'hd0 : c[0:7] = 8'h67;
			8'hd1 : c[0:7] = 8'h6a;
			8'hd2 : c[0:7] = 8'h7d;
			8'hd3 : c[0:7] = 8'h70;
			8'hd4 : c[0:7] = 8'h53;
			8'hd5 : c[0:7] = 8'h5e;
			8'hd6 : c[0:7] = 8'h49;
			8'hd7 : c[0:7] = 8'h44;
			8'hd8 : c[0:7] = 8'hf;
			8'hd9 : c[0:7] = 8'h2;
			8'hda : c[0:7] = 8'h15;
			8'hdb : c[0:7] = 8'h18;
			8'hdc : c[0:7] = 8'h3b;
			8'hdd : c[0:7] = 8'h36;
			8'hde : c[0:7] = 8'h21;
			8'hdf : c[0:7] = 8'h2c;
			8'he0 : c[0:7] = 8'hc;
			8'he1 : c[0:7] = 8'h1;
			8'he2 : c[0:7] = 8'h16;
			8'he3 : c[0:7] = 8'h1b;
			8'he4 : c[0:7] = 8'h38;
			8'he5 : c[0:7] = 8'h35;
			8'he6 : c[0:7] = 8'h22;
			8'he7 : c[0:7] = 8'h2f;
			8'he8 : c[0:7] = 8'h64;
			8'he9 : c[0:7] = 8'h69;
			8'hea : c[0:7] = 8'h7e;
			8'heb : c[0:7] = 8'h73;
			8'hec : c[0:7] = 8'h50;
			8'hed : c[0:7] = 8'h5d;
			8'hee : c[0:7] = 8'h4a;
			8'hef : c[0:7] = 8'h47;
			8'hf0 : c[0:7] = 8'hdc;
			8'hf1 : c[0:7] = 8'hd1;
			8'hf2 : c[0:7] = 8'hc6;
			8'hf3 : c[0:7] = 8'hcb;
			8'hf4 : c[0:7] = 8'he8;
			8'hf5 : c[0:7] = 8'he5;
			8'hf6 : c[0:7] = 8'hf2;
			8'hf7 : c[0:7] = 8'hff;
			8'hf8 : c[0:7] = 8'hb4;
			8'hf9 : c[0:7] = 8'hb9;
			8'hfa : c[0:7] = 8'hae;
			8'hfb : c[0:7] = 8'ha3;
			8'hfc : c[0:7] = 8'h80;
			8'hfd : c[0:7] = 8'h8d;
			8'hfe : c[0:7] = 8'h9a;
			8'hff : c[0:7] = 8'h97;			
        endcase
    end

    assign output_row = a ^ b ^ c ^ d;
    
endmodule


module MixColumn3RowInverse (
    input wire [0:31] row,
    output wire [0:7] output_row
);
    reg [0:7] a, b, c, d;

    // Multiplication with 13
    always @(row[0:7]) begin
        case (row[0:7])
            			8'h0 : c[0:7] = 8'h0;
			8'h1 : c[0:7] = 8'hd;
			8'h2 : c[0:7] = 8'h1a;
			8'h3 : c[0:7] = 8'h17;
			8'h4 : c[0:7] = 8'h34;
			8'h5 : c[0:7] = 8'h39;
			8'h6 : c[0:7] = 8'h2e;
			8'h7 : c[0:7] = 8'h23;
			8'h8 : c[0:7] = 8'h68;
			8'h9 : c[0:7] = 8'h65;
			8'ha : c[0:7] = 8'h72;
			8'hb : c[0:7] = 8'h7f;
			8'hc : c[0:7] = 8'h5c;
			8'hd : c[0:7] = 8'h51;
			8'he : c[0:7] = 8'h46;
			8'hf : c[0:7] = 8'h4b;
			8'h10 : c[0:7] = 8'hd0;
			8'h11 : c[0:7] = 8'hdd;
			8'h12 : c[0:7] = 8'hca;
			8'h13 : c[0:7] = 8'hc7;
			8'h14 : c[0:7] = 8'he4;
			8'h15 : c[0:7] = 8'he9;
			8'h16 : c[0:7] = 8'hfe;
			8'h17 : c[0:7] = 8'hf3;
			8'h18 : c[0:7] = 8'hb8;
			8'h19 : c[0:7] = 8'hb5;
			8'h1a : c[0:7] = 8'ha2;
			8'h1b : c[0:7] = 8'haf;
			8'h1c : c[0:7] = 8'h8c;
			8'h1d : c[0:7] = 8'h81;
			8'h1e : c[0:7] = 8'h96;
			8'h1f : c[0:7] = 8'h9b;
			8'h20 : c[0:7] = 8'hbb;
			8'h21 : c[0:7] = 8'hb6;
			8'h22 : c[0:7] = 8'ha1;
			8'h23 : c[0:7] = 8'hac;
			8'h24 : c[0:7] = 8'h8f;
			8'h25 : c[0:7] = 8'h82;
			8'h26 : c[0:7] = 8'h95;
			8'h27 : c[0:7] = 8'h98;
			8'h28 : c[0:7] = 8'hd3;
			8'h29 : c[0:7] = 8'hde;
			8'h2a : c[0:7] = 8'hc9;
			8'h2b : c[0:7] = 8'hc4;
			8'h2c : c[0:7] = 8'he7;
			8'h2d : c[0:7] = 8'hea;
			8'h2e : c[0:7] = 8'hfd;
			8'h2f : c[0:7] = 8'hf0;
			8'h30 : c[0:7] = 8'h6b;
			8'h31 : c[0:7] = 8'h66;
			8'h32 : c[0:7] = 8'h71;
			8'h33 : c[0:7] = 8'h7c;
			8'h34 : c[0:7] = 8'h5f;
			8'h35 : c[0:7] = 8'h52;
			8'h36 : c[0:7] = 8'h45;
			8'h37 : c[0:7] = 8'h48;
			8'h38 : c[0:7] = 8'h3;
			8'h39 : c[0:7] = 8'he;
			8'h3a : c[0:7] = 8'h19;
			8'h3b : c[0:7] = 8'h14;
			8'h3c : c[0:7] = 8'h37;
			8'h3d : c[0:7] = 8'h3a;
			8'h3e : c[0:7] = 8'h2d;
			8'h3f : c[0:7] = 8'h20;
			8'h40 : c[0:7] = 8'h6d;
			8'h41 : c[0:7] = 8'h60;
			8'h42 : c[0:7] = 8'h77;
			8'h43 : c[0:7] = 8'h7a;
			8'h44 : c[0:7] = 8'h59;
			8'h45 : c[0:7] = 8'h54;
			8'h46 : c[0:7] = 8'h43;
			8'h47 : c[0:7] = 8'h4e;
			8'h48 : c[0:7] = 8'h5;
			8'h49 : c[0:7] = 8'h8;
			8'h4a : c[0:7] = 8'h1f;
			8'h4b : c[0:7] = 8'h12;
			8'h4c : c[0:7] = 8'h31;
			8'h4d : c[0:7] = 8'h3c;
			8'h4e : c[0:7] = 8'h2b;
			8'h4f : c[0:7] = 8'h26;
			8'h50 : c[0:7] = 8'hbd;
			8'h51 : c[0:7] = 8'hb0;
			8'h52 : c[0:7] = 8'ha7;
			8'h53 : c[0:7] = 8'haa;
			8'h54 : c[0:7] = 8'h89;
			8'h55 : c[0:7] = 8'h84;
			8'h56 : c[0:7] = 8'h93;
			8'h57 : c[0:7] = 8'h9e;
			8'h58 : c[0:7] = 8'hd5;
			8'h59 : c[0:7] = 8'hd8;
			8'h5a : c[0:7] = 8'hcf;
			8'h5b : c[0:7] = 8'hc2;
			8'h5c : c[0:7] = 8'he1;
			8'h5d : c[0:7] = 8'hec;
			8'h5e : c[0:7] = 8'hfb;
			8'h5f : c[0:7] = 8'hf6;
			8'h60 : c[0:7] = 8'hd6;
			8'h61 : c[0:7] = 8'hdb;
			8'h62 : c[0:7] = 8'hcc;
			8'h63 : c[0:7] = 8'hc1;
			8'h64 : c[0:7] = 8'he2;
			8'h65 : c[0:7] = 8'hef;
			8'h66 : c[0:7] = 8'hf8;
			8'h67 : c[0:7] = 8'hf5;
			8'h68 : c[0:7] = 8'hbe;
			8'h69 : c[0:7] = 8'hb3;
			8'h6a : c[0:7] = 8'ha4;
			8'h6b : c[0:7] = 8'ha9;
			8'h6c : c[0:7] = 8'h8a;
			8'h6d : c[0:7] = 8'h87;
			8'h6e : c[0:7] = 8'h90;
			8'h6f : c[0:7] = 8'h9d;
			8'h70 : c[0:7] = 8'h6;
			8'h71 : c[0:7] = 8'hb;
			8'h72 : c[0:7] = 8'h1c;
			8'h73 : c[0:7] = 8'h11;
			8'h74 : c[0:7] = 8'h32;
			8'h75 : c[0:7] = 8'h3f;
			8'h76 : c[0:7] = 8'h28;
			8'h77 : c[0:7] = 8'h25;
			8'h78 : c[0:7] = 8'h6e;
			8'h79 : c[0:7] = 8'h63;
			8'h7a : c[0:7] = 8'h74;
			8'h7b : c[0:7] = 8'h79;
			8'h7c : c[0:7] = 8'h5a;
			8'h7d : c[0:7] = 8'h57;
			8'h7e : c[0:7] = 8'h40;
			8'h7f : c[0:7] = 8'h4d;
			8'h80 : c[0:7] = 8'hda;
			8'h81 : c[0:7] = 8'hd7;
			8'h82 : c[0:7] = 8'hc0;
			8'h83 : c[0:7] = 8'hcd;
			8'h84 : c[0:7] = 8'hee;
			8'h85 : c[0:7] = 8'he3;
			8'h86 : c[0:7] = 8'hf4;
			8'h87 : c[0:7] = 8'hf9;
			8'h88 : c[0:7] = 8'hb2;
			8'h89 : c[0:7] = 8'hbf;
			8'h8a : c[0:7] = 8'ha8;
			8'h8b : c[0:7] = 8'ha5;
			8'h8c : c[0:7] = 8'h86;
			8'h8d : c[0:7] = 8'h8b;
			8'h8e : c[0:7] = 8'h9c;
			8'h8f : c[0:7] = 8'h91;
			8'h90 : c[0:7] = 8'ha;
			8'h91 : c[0:7] = 8'h7;
			8'h92 : c[0:7] = 8'h10;
			8'h93 : c[0:7] = 8'h1d;
			8'h94 : c[0:7] = 8'h3e;
			8'h95 : c[0:7] = 8'h33;
			8'h96 : c[0:7] = 8'h24;
			8'h97 : c[0:7] = 8'h29;
			8'h98 : c[0:7] = 8'h62;
			8'h99 : c[0:7] = 8'h6f;
			8'h9a : c[0:7] = 8'h78;
			8'h9b : c[0:7] = 8'h75;
			8'h9c : c[0:7] = 8'h56;
			8'h9d : c[0:7] = 8'h5b;
			8'h9e : c[0:7] = 8'h4c;
			8'h9f : c[0:7] = 8'h41;
			8'ha0 : c[0:7] = 8'h61;
			8'ha1 : c[0:7] = 8'h6c;
			8'ha2 : c[0:7] = 8'h7b;
			8'ha3 : c[0:7] = 8'h76;
			8'ha4 : c[0:7] = 8'h55;
			8'ha5 : c[0:7] = 8'h58;
			8'ha6 : c[0:7] = 8'h4f;
			8'ha7 : c[0:7] = 8'h42;
			8'ha8 : c[0:7] = 8'h9;
			8'ha9 : c[0:7] = 8'h4;
			8'haa : c[0:7] = 8'h13;
			8'hab : c[0:7] = 8'h1e;
			8'hac : c[0:7] = 8'h3d;
			8'had : c[0:7] = 8'h30;
			8'hae : c[0:7] = 8'h27;
			8'haf : c[0:7] = 8'h2a;
			8'hb0 : c[0:7] = 8'hb1;
			8'hb1 : c[0:7] = 8'hbc;
			8'hb2 : c[0:7] = 8'hab;
			8'hb3 : c[0:7] = 8'ha6;
			8'hb4 : c[0:7] = 8'h85;
			8'hb5 : c[0:7] = 8'h88;
			8'hb6 : c[0:7] = 8'h9f;
			8'hb7 : c[0:7] = 8'h92;
			8'hb8 : c[0:7] = 8'hd9;
			8'hb9 : c[0:7] = 8'hd4;
			8'hba : c[0:7] = 8'hc3;
			8'hbb : c[0:7] = 8'hce;
			8'hbc : c[0:7] = 8'hed;
			8'hbd : c[0:7] = 8'he0;
			8'hbe : c[0:7] = 8'hf7;
			8'hbf : c[0:7] = 8'hfa;
			8'hc0 : c[0:7] = 8'hb7;
			8'hc1 : c[0:7] = 8'hba;
			8'hc2 : c[0:7] = 8'had;
			8'hc3 : c[0:7] = 8'ha0;
			8'hc4 : c[0:7] = 8'h83;
			8'hc5 : c[0:7] = 8'h8e;
			8'hc6 : c[0:7] = 8'h99;
			8'hc7 : c[0:7] = 8'h94;
			8'hc8 : c[0:7] = 8'hdf;
			8'hc9 : c[0:7] = 8'hd2;
			8'hca : c[0:7] = 8'hc5;
			8'hcb : c[0:7] = 8'hc8;
			8'hcc : c[0:7] = 8'heb;
			8'hcd : c[0:7] = 8'he6;
			8'hce : c[0:7] = 8'hf1;
			8'hcf : c[0:7] = 8'hfc;
			8'hd0 : c[0:7] = 8'h67;
			8'hd1 : c[0:7] = 8'h6a;
			8'hd2 : c[0:7] = 8'h7d;
			8'hd3 : c[0:7] = 8'h70;
			8'hd4 : c[0:7] = 8'h53;
			8'hd5 : c[0:7] = 8'h5e;
			8'hd6 : c[0:7] = 8'h49;
			8'hd7 : c[0:7] = 8'h44;
			8'hd8 : c[0:7] = 8'hf;
			8'hd9 : c[0:7] = 8'h2;
			8'hda : c[0:7] = 8'h15;
			8'hdb : c[0:7] = 8'h18;
			8'hdc : c[0:7] = 8'h3b;
			8'hdd : c[0:7] = 8'h36;
			8'hde : c[0:7] = 8'h21;
			8'hdf : c[0:7] = 8'h2c;
			8'he0 : c[0:7] = 8'hc;
			8'he1 : c[0:7] = 8'h1;
			8'he2 : c[0:7] = 8'h16;
			8'he3 : c[0:7] = 8'h1b;
			8'he4 : c[0:7] = 8'h38;
			8'he5 : c[0:7] = 8'h35;
			8'he6 : c[0:7] = 8'h22;
			8'he7 : c[0:7] = 8'h2f;
			8'he8 : c[0:7] = 8'h64;
			8'he9 : c[0:7] = 8'h69;
			8'hea : c[0:7] = 8'h7e;
			8'heb : c[0:7] = 8'h73;
			8'hec : c[0:7] = 8'h50;
			8'hed : c[0:7] = 8'h5d;
			8'hee : c[0:7] = 8'h4a;
			8'hef : c[0:7] = 8'h47;
			8'hf0 : c[0:7] = 8'hdc;
			8'hf1 : c[0:7] = 8'hd1;
			8'hf2 : c[0:7] = 8'hc6;
			8'hf3 : c[0:7] = 8'hcb;
			8'hf4 : c[0:7] = 8'he8;
			8'hf5 : c[0:7] = 8'he5;
			8'hf6 : c[0:7] = 8'hf2;
			8'hf7 : c[0:7] = 8'hff;
			8'hf8 : c[0:7] = 8'hb4;
			8'hf9 : c[0:7] = 8'hb9;
			8'hfa : c[0:7] = 8'hae;
			8'hfb : c[0:7] = 8'ha3;
			8'hfc : c[0:7] = 8'h80;
			8'hfd : c[0:7] = 8'h8d;
			8'hfe : c[0:7] = 8'h9a;
			8'hff : c[0:7] = 8'h97;
        endcase
    end

    // Multiplication with 9
    always @(row[8:15]) begin
        case (row[8:15])
            8'h0 : d[0:7] = 8'h0;
			8'h1 : d[0:7] = 8'h9;
			8'h2 : d[0:7] = 8'h12;
			8'h3 : d[0:7] = 8'h1b;
			8'h4 : d[0:7] = 8'h24;
			8'h5 : d[0:7] = 8'h2d;
			8'h6 : d[0:7] = 8'h36;
			8'h7 : d[0:7] = 8'h3f;
			8'h8 : d[0:7] = 8'h48;
			8'h9 : d[0:7] = 8'h41;
			8'ha : d[0:7] = 8'h5a;
			8'hb : d[0:7] = 8'h53;
			8'hc : d[0:7] = 8'h6c;
			8'hd : d[0:7] = 8'h65;
			8'he : d[0:7] = 8'h7e;
			8'hf : d[0:7] = 8'h77;
			8'h10 : d[0:7] = 8'h90;
			8'h11 : d[0:7] = 8'h99;
			8'h12 : d[0:7] = 8'h82;
			8'h13 : d[0:7] = 8'h8b;
			8'h14 : d[0:7] = 8'hb4;
			8'h15 : d[0:7] = 8'hbd;
			8'h16 : d[0:7] = 8'ha6;
			8'h17 : d[0:7] = 8'haf;
			8'h18 : d[0:7] = 8'hd8;
			8'h19 : d[0:7] = 8'hd1;
			8'h1a : d[0:7] = 8'hca;
			8'h1b : d[0:7] = 8'hc3;
			8'h1c : d[0:7] = 8'hfc;
			8'h1d : d[0:7] = 8'hf5;
			8'h1e : d[0:7] = 8'hee;
			8'h1f : d[0:7] = 8'he7;
			8'h20 : d[0:7] = 8'h3b;
			8'h21 : d[0:7] = 8'h32;
			8'h22 : d[0:7] = 8'h29;
			8'h23 : d[0:7] = 8'h20;
			8'h24 : d[0:7] = 8'h1f;
			8'h25 : d[0:7] = 8'h16;
			8'h26 : d[0:7] = 8'hd;
			8'h27 : d[0:7] = 8'h4;
			8'h28 : d[0:7] = 8'h73;
			8'h29 : d[0:7] = 8'h7a;
			8'h2a : d[0:7] = 8'h61;
			8'h2b : d[0:7] = 8'h68;
			8'h2c : d[0:7] = 8'h57;
			8'h2d : d[0:7] = 8'h5e;
			8'h2e : d[0:7] = 8'h45;
			8'h2f : d[0:7] = 8'h4c;
			8'h30 : d[0:7] = 8'hab;
			8'h31 : d[0:7] = 8'ha2;
			8'h32 : d[0:7] = 8'hb9;
			8'h33 : d[0:7] = 8'hb0;
			8'h34 : d[0:7] = 8'h8f;
			8'h35 : d[0:7] = 8'h86;
			8'h36 : d[0:7] = 8'h9d;
			8'h37 : d[0:7] = 8'h94;
			8'h38 : d[0:7] = 8'he3;
			8'h39 : d[0:7] = 8'hea;
			8'h3a : d[0:7] = 8'hf1;
			8'h3b : d[0:7] = 8'hf8;
			8'h3c : d[0:7] = 8'hc7;
			8'h3d : d[0:7] = 8'hce;
			8'h3e : d[0:7] = 8'hd5;
			8'h3f : d[0:7] = 8'hdc;
			8'h40 : d[0:7] = 8'h76;
			8'h41 : d[0:7] = 8'h7f;
			8'h42 : d[0:7] = 8'h64;
			8'h43 : d[0:7] = 8'h6d;
			8'h44 : d[0:7] = 8'h52;
			8'h45 : d[0:7] = 8'h5b;
			8'h46 : d[0:7] = 8'h40;
			8'h47 : d[0:7] = 8'h49;
			8'h48 : d[0:7] = 8'h3e;
			8'h49 : d[0:7] = 8'h37;
			8'h4a : d[0:7] = 8'h2c;
			8'h4b : d[0:7] = 8'h25;
			8'h4c : d[0:7] = 8'h1a;
			8'h4d : d[0:7] = 8'h13;
			8'h4e : d[0:7] = 8'h8;
			8'h4f : d[0:7] = 8'h1;
			8'h50 : d[0:7] = 8'he6;
			8'h51 : d[0:7] = 8'hef;
			8'h52 : d[0:7] = 8'hf4;
			8'h53 : d[0:7] = 8'hfd;
			8'h54 : d[0:7] = 8'hc2;
			8'h55 : d[0:7] = 8'hcb;
			8'h56 : d[0:7] = 8'hd0;
			8'h57 : d[0:7] = 8'hd9;
			8'h58 : d[0:7] = 8'hae;
			8'h59 : d[0:7] = 8'ha7;
			8'h5a : d[0:7] = 8'hbc;
			8'h5b : d[0:7] = 8'hb5;
			8'h5c : d[0:7] = 8'h8a;
			8'h5d : d[0:7] = 8'h83;
			8'h5e : d[0:7] = 8'h98;
			8'h5f : d[0:7] = 8'h91;
			8'h60 : d[0:7] = 8'h4d;
			8'h61 : d[0:7] = 8'h44;
			8'h62 : d[0:7] = 8'h5f;
			8'h63 : d[0:7] = 8'h56;
			8'h64 : d[0:7] = 8'h69;
			8'h65 : d[0:7] = 8'h60;
			8'h66 : d[0:7] = 8'h7b;
			8'h67 : d[0:7] = 8'h72;
			8'h68 : d[0:7] = 8'h5;
			8'h69 : d[0:7] = 8'hc;
			8'h6a : d[0:7] = 8'h17;
			8'h6b : d[0:7] = 8'h1e;
			8'h6c : d[0:7] = 8'h21;
			8'h6d : d[0:7] = 8'h28;
			8'h6e : d[0:7] = 8'h33;
			8'h6f : d[0:7] = 8'h3a;
			8'h70 : d[0:7] = 8'hdd;
			8'h71 : d[0:7] = 8'hd4;
			8'h72 : d[0:7] = 8'hcf;
			8'h73 : d[0:7] = 8'hc6;
			8'h74 : d[0:7] = 8'hf9;
			8'h75 : d[0:7] = 8'hf0;
			8'h76 : d[0:7] = 8'heb;
			8'h77 : d[0:7] = 8'he2;
			8'h78 : d[0:7] = 8'h95;
			8'h79 : d[0:7] = 8'h9c;
			8'h7a : d[0:7] = 8'h87;
			8'h7b : d[0:7] = 8'h8e;
			8'h7c : d[0:7] = 8'hb1;
			8'h7d : d[0:7] = 8'hb8;
			8'h7e : d[0:7] = 8'ha3;
			8'h7f : d[0:7] = 8'haa;
			8'h80 : d[0:7] = 8'hec;
			8'h81 : d[0:7] = 8'he5;
			8'h82 : d[0:7] = 8'hfe;
			8'h83 : d[0:7] = 8'hf7;
			8'h84 : d[0:7] = 8'hc8;
			8'h85 : d[0:7] = 8'hc1;
			8'h86 : d[0:7] = 8'hda;
			8'h87 : d[0:7] = 8'hd3;
			8'h88 : d[0:7] = 8'ha4;
			8'h89 : d[0:7] = 8'had;
			8'h8a : d[0:7] = 8'hb6;
			8'h8b : d[0:7] = 8'hbf;
			8'h8c : d[0:7] = 8'h80;
			8'h8d : d[0:7] = 8'h89;
			8'h8e : d[0:7] = 8'h92;
			8'h8f : d[0:7] = 8'h9b;
			8'h90 : d[0:7] = 8'h7c;
			8'h91 : d[0:7] = 8'h75;
			8'h92 : d[0:7] = 8'h6e;
			8'h93 : d[0:7] = 8'h67;
			8'h94 : d[0:7] = 8'h58;
			8'h95 : d[0:7] = 8'h51;
			8'h96 : d[0:7] = 8'h4a;
			8'h97 : d[0:7] = 8'h43;
			8'h98 : d[0:7] = 8'h34;
			8'h99 : d[0:7] = 8'h3d;
			8'h9a : d[0:7] = 8'h26;
			8'h9b : d[0:7] = 8'h2f;
			8'h9c : d[0:7] = 8'h10;
			8'h9d : d[0:7] = 8'h19;
			8'h9e : d[0:7] = 8'h2;
			8'h9f : d[0:7] = 8'hb;
			8'ha0 : d[0:7] = 8'hd7;
			8'ha1 : d[0:7] = 8'hde;
			8'ha2 : d[0:7] = 8'hc5;
			8'ha3 : d[0:7] = 8'hcc;
			8'ha4 : d[0:7] = 8'hf3;
			8'ha5 : d[0:7] = 8'hfa;
			8'ha6 : d[0:7] = 8'he1;
			8'ha7 : d[0:7] = 8'he8;
			8'ha8 : d[0:7] = 8'h9f;
			8'ha9 : d[0:7] = 8'h96;
			8'haa : d[0:7] = 8'h8d;
			8'hab : d[0:7] = 8'h84;
			8'hac : d[0:7] = 8'hbb;
			8'had : d[0:7] = 8'hb2;
			8'hae : d[0:7] = 8'ha9;
			8'haf : d[0:7] = 8'ha0;
			8'hb0 : d[0:7] = 8'h47;
			8'hb1 : d[0:7] = 8'h4e;
			8'hb2 : d[0:7] = 8'h55;
			8'hb3 : d[0:7] = 8'h5c;
			8'hb4 : d[0:7] = 8'h63;
			8'hb5 : d[0:7] = 8'h6a;
			8'hb6 : d[0:7] = 8'h71;
			8'hb7 : d[0:7] = 8'h78;
			8'hb8 : d[0:7] = 8'hf;
			8'hb9 : d[0:7] = 8'h6;
			8'hba : d[0:7] = 8'h1d;
			8'hbb : d[0:7] = 8'h14;
			8'hbc : d[0:7] = 8'h2b;
			8'hbd : d[0:7] = 8'h22;
			8'hbe : d[0:7] = 8'h39;
			8'hbf : d[0:7] = 8'h30;
			8'hc0 : d[0:7] = 8'h9a;
			8'hc1 : d[0:7] = 8'h93;
			8'hc2 : d[0:7] = 8'h88;
			8'hc3 : d[0:7] = 8'h81;
			8'hc4 : d[0:7] = 8'hbe;
			8'hc5 : d[0:7] = 8'hb7;
			8'hc6 : d[0:7] = 8'hac;
			8'hc7 : d[0:7] = 8'ha5;
			8'hc8 : d[0:7] = 8'hd2;
			8'hc9 : d[0:7] = 8'hdb;
			8'hca : d[0:7] = 8'hc0;
			8'hcb : d[0:7] = 8'hc9;
			8'hcc : d[0:7] = 8'hf6;
			8'hcd : d[0:7] = 8'hff;
			8'hce : d[0:7] = 8'he4;
			8'hcf : d[0:7] = 8'hed;
			8'hd0 : d[0:7] = 8'ha;
			8'hd1 : d[0:7] = 8'h3;
			8'hd2 : d[0:7] = 8'h18;
			8'hd3 : d[0:7] = 8'h11;
			8'hd4 : d[0:7] = 8'h2e;
			8'hd5 : d[0:7] = 8'h27;
			8'hd6 : d[0:7] = 8'h3c;
			8'hd7 : d[0:7] = 8'h35;
			8'hd8 : d[0:7] = 8'h42;
			8'hd9 : d[0:7] = 8'h4b;
			8'hda : d[0:7] = 8'h50;
			8'hdb : d[0:7] = 8'h59;
			8'hdc : d[0:7] = 8'h66;
			8'hdd : d[0:7] = 8'h6f;
			8'hde : d[0:7] = 8'h74;
			8'hdf : d[0:7] = 8'h7d;
			8'he0 : d[0:7] = 8'ha1;
			8'he1 : d[0:7] = 8'ha8;
			8'he2 : d[0:7] = 8'hb3;
			8'he3 : d[0:7] = 8'hba;
			8'he4 : d[0:7] = 8'h85;
			8'he5 : d[0:7] = 8'h8c;
			8'he6 : d[0:7] = 8'h97;
			8'he7 : d[0:7] = 8'h9e;
			8'he8 : d[0:7] = 8'he9;
			8'he9 : d[0:7] = 8'he0;
			8'hea : d[0:7] = 8'hfb;
			8'heb : d[0:7] = 8'hf2;
			8'hec : d[0:7] = 8'hcd;
			8'hed : d[0:7] = 8'hc4;
			8'hee : d[0:7] = 8'hdf;
			8'hef : d[0:7] = 8'hd6;
			8'hf0 : d[0:7] = 8'h31;
			8'hf1 : d[0:7] = 8'h38;
			8'hf2 : d[0:7] = 8'h23;
			8'hf3 : d[0:7] = 8'h2a;
			8'hf4 : d[0:7] = 8'h15;
			8'hf5 : d[0:7] = 8'h1c;
			8'hf6 : d[0:7] = 8'h7;
			8'hf7 : d[0:7] = 8'he;
			8'hf8 : d[0:7] = 8'h79;
			8'hf9 : d[0:7] = 8'h70;
			8'hfa : d[0:7] = 8'h6b;
			8'hfb : d[0:7] = 8'h62;
			8'hfc : d[0:7] = 8'h5d;
			8'hfd : d[0:7] = 8'h54;
			8'hfe : d[0:7] = 8'h4f;
			8'hff : d[0:7] = 8'h46;
        endcase
    end

    // Multiplication with 14
    always @(row[16:23]) begin
        case (row[16:23])
			            8'h0 : a[0:7] = 8'h0;
            8'h1 : a[0:7] = 8'he;
            8'h2 : a[0:7] = 8'h1c;
            8'h3 : a[0:7] = 8'h12;
            8'h4 : a[0:7] = 8'h38;
            8'h5 : a[0:7] = 8'h36;
            8'h6 : a[0:7] = 8'h24;
            8'h7 : a[0:7] = 8'h2a;
            8'h8 : a[0:7] = 8'h70;
            8'h9 : a[0:7] = 8'h7e;
            8'ha : a[0:7] = 8'h6c;
            8'hb : a[0:7] = 8'h62;
            8'hc : a[0:7] = 8'h48;
            8'hd : a[0:7] = 8'h46;
            8'he : a[0:7] = 8'h54;
            8'hf : a[0:7] = 8'h5a;
            8'h10 : a[0:7] = 8'he0;
            8'h11 : a[0:7] = 8'hee;
            8'h12 : a[0:7] = 8'hfc;
            8'h13 : a[0:7] = 8'hf2;
            8'h14 : a[0:7] = 8'hd8;
            8'h15 : a[0:7] = 8'hd6;
            8'h16 : a[0:7] = 8'hc4;
            8'h17 : a[0:7] = 8'hca;
            8'h18 : a[0:7] = 8'h90;
            8'h19 : a[0:7] = 8'h9e;
            8'h1a : a[0:7] = 8'h8c;
            8'h1b : a[0:7] = 8'h82;
            8'h1c : a[0:7] = 8'ha8;
            8'h1d : a[0:7] = 8'ha6;
            8'h1e : a[0:7] = 8'hb4;
            8'h1f : a[0:7] = 8'hba;
            8'h20 : a[0:7] = 8'hdb;
            8'h21 : a[0:7] = 8'hd5;
            8'h22 : a[0:7] = 8'hc7;
            8'h23 : a[0:7] = 8'hc9;
            8'h24 : a[0:7] = 8'he3;
            8'h25 : a[0:7] = 8'hed;
            8'h26 : a[0:7] = 8'hff;
            8'h27 : a[0:7] = 8'hf1;
            8'h28 : a[0:7] = 8'hab;
            8'h29 : a[0:7] = 8'ha5;
            8'h2a : a[0:7] = 8'hb7;
            8'h2b : a[0:7] = 8'hb9;
            8'h2c : a[0:7] = 8'h93;
            8'h2d : a[0:7] = 8'h9d;
            8'h2e : a[0:7] = 8'h8f;
            8'h2f : a[0:7] = 8'h81;
            8'h30 : a[0:7] = 8'h3b;
            8'h31 : a[0:7] = 8'h35;
            8'h32 : a[0:7] = 8'h27;
            8'h33 : a[0:7] = 8'h29;
            8'h34 : a[0:7] = 8'h3;
            8'h35 : a[0:7] = 8'hd;
            8'h36 : a[0:7] = 8'h1f;
            8'h37 : a[0:7] = 8'h11;
            8'h38 : a[0:7] = 8'h4b;
            8'h39 : a[0:7] = 8'h45;
            8'h3a : a[0:7] = 8'h57;
            8'h3b : a[0:7] = 8'h59;
            8'h3c : a[0:7] = 8'h73;
            8'h3d : a[0:7] = 8'h7d;
            8'h3e : a[0:7] = 8'h6f;
            8'h3f : a[0:7] = 8'h61;
            8'h40 : a[0:7] = 8'had;
            8'h41 : a[0:7] = 8'ha3;
            8'h42 : a[0:7] = 8'hb1;
            8'h43 : a[0:7] = 8'hbf;
            8'h44 : a[0:7] = 8'h95;
            8'h45 : a[0:7] = 8'h9b;
            8'h46 : a[0:7] = 8'h89;
            8'h47 : a[0:7] = 8'h87;
            8'h48 : a[0:7] = 8'hdd;
            8'h49 : a[0:7] = 8'hd3;
            8'h4a : a[0:7] = 8'hc1;
            8'h4b : a[0:7] = 8'hcf;
            8'h4c : a[0:7] = 8'he5;
            8'h4d : a[0:7] = 8'heb;
            8'h4e : a[0:7] = 8'hf9;
            8'h4f : a[0:7] = 8'hf7;
            8'h50 : a[0:7] = 8'h4d;
            8'h51 : a[0:7] = 8'h43;
            8'h52 : a[0:7] = 8'h51;
            8'h53 : a[0:7] = 8'h5f;
            8'h54 : a[0:7] = 8'h75;
            8'h55 : a[0:7] = 8'h7b;
            8'h56 : a[0:7] = 8'h69;
            8'h57 : a[0:7] = 8'h67;
            8'h58 : a[0:7] = 8'h3d;
            8'h59 : a[0:7] = 8'h33;
            8'h5a : a[0:7] = 8'h21;
            8'h5b : a[0:7] = 8'h2f;
            8'h5c : a[0:7] = 8'h5;
            8'h5d : a[0:7] = 8'hb;
            8'h5e : a[0:7] = 8'h19;
            8'h5f : a[0:7] = 8'h17;
            8'h60 : a[0:7] = 8'h76;
            8'h61 : a[0:7] = 8'h78;
            8'h62 : a[0:7] = 8'h6a;
            8'h63 : a[0:7] = 8'h64;
            8'h64 : a[0:7] = 8'h4e;
            8'h65 : a[0:7] = 8'h40;
            8'h66 : a[0:7] = 8'h52;
            8'h67 : a[0:7] = 8'h5c;
            8'h68 : a[0:7] = 8'h6;
            8'h69 : a[0:7] = 8'h8;
            8'h6a : a[0:7] = 8'h1a;
            8'h6b : a[0:7] = 8'h14;
            8'h6c : a[0:7] = 8'h3e;
            8'h6d : a[0:7] = 8'h30;
            8'h6e : a[0:7] = 8'h22;
            8'h6f : a[0:7] = 8'h2c;
            8'h70 : a[0:7] = 8'h96;
            8'h71 : a[0:7] = 8'h98;
            8'h72 : a[0:7] = 8'h8a;
            8'h73 : a[0:7] = 8'h84;
            8'h74 : a[0:7] = 8'hae;
            8'h75 : a[0:7] = 8'ha0;
            8'h76 : a[0:7] = 8'hb2;
            8'h77 : a[0:7] = 8'hbc;
            8'h78 : a[0:7] = 8'he6;
            8'h79 : a[0:7] = 8'he8;
            8'h7a : a[0:7] = 8'hfa;
            8'h7b : a[0:7] = 8'hf4;
            8'h7c : a[0:7] = 8'hde;
            8'h7d : a[0:7] = 8'hd0;
            8'h7e : a[0:7] = 8'hc2;
            8'h7f : a[0:7] = 8'hcc;
            8'h80 : a[0:7] = 8'h41;
            8'h81 : a[0:7] = 8'h4f;
            8'h82 : a[0:7] = 8'h5d;
            8'h83 : a[0:7] = 8'h53;
            8'h84 : a[0:7] = 8'h79;
            8'h85 : a[0:7] = 8'h77;
            8'h86 : a[0:7] = 8'h65;
            8'h87 : a[0:7] = 8'h6b;
            8'h88 : a[0:7] = 8'h31;
            8'h89 : a[0:7] = 8'h3f;
            8'h8a : a[0:7] = 8'h2d;
            8'h8b : a[0:7] = 8'h23;
            8'h8c : a[0:7] = 8'h9;
            8'h8d : a[0:7] = 8'h7;
            8'h8e : a[0:7] = 8'h15;
            8'h8f : a[0:7] = 8'h1b;
            8'h90 : a[0:7] = 8'ha1;
            8'h91 : a[0:7] = 8'haf;
            8'h92 : a[0:7] = 8'hbd;
            8'h93 : a[0:7] = 8'hb3;
            8'h94 : a[0:7] = 8'h99;
            8'h95 : a[0:7] = 8'h97;
            8'h96 : a[0:7] = 8'h85;
            8'h97 : a[0:7] = 8'h8b;
            8'h98 : a[0:7] = 8'hd1;
            8'h99 : a[0:7] = 8'hdf;
            8'h9a : a[0:7] = 8'hcd;
            8'h9b : a[0:7] = 8'hc3;
            8'h9c : a[0:7] = 8'he9;
            8'h9d : a[0:7] = 8'he7;
            8'h9e : a[0:7] = 8'hf5;
            8'h9f : a[0:7] = 8'hfb;
            8'ha0 : a[0:7] = 8'h9a;
            8'ha1 : a[0:7] = 8'h94;
            8'ha2 : a[0:7] = 8'h86;
            8'ha3 : a[0:7] = 8'h88;
            8'ha4 : a[0:7] = 8'ha2;
            8'ha5 : a[0:7] = 8'hac;
            8'ha6 : a[0:7] = 8'hbe;
            8'ha7 : a[0:7] = 8'hb0;
            8'ha8 : a[0:7] = 8'hea;
            8'ha9 : a[0:7] = 8'he4;
            8'haa : a[0:7] = 8'hf6;
            8'hab : a[0:7] = 8'hf8;
            8'hac : a[0:7] = 8'hd2;
            8'had : a[0:7] = 8'hdc;
            8'hae : a[0:7] = 8'hce;
            8'haf : a[0:7] = 8'hc0;
            8'hb0 : a[0:7] = 8'h7a;
            8'hb1 : a[0:7] = 8'h74;
            8'hb2 : a[0:7] = 8'h66;
            8'hb3 : a[0:7] = 8'h68;
            8'hb4 : a[0:7] = 8'h42;
            8'hb5 : a[0:7] = 8'h4c;
            8'hb6 : a[0:7] = 8'h5e;
            8'hb7 : a[0:7] = 8'h50;
            8'hb8 : a[0:7] = 8'ha;
            8'hb9 : a[0:7] = 8'h4;
            8'hba : a[0:7] = 8'h16;
            8'hbb : a[0:7] = 8'h18;
            8'hbc : a[0:7] = 8'h32;
            8'hbd : a[0:7] = 8'h3c;
            8'hbe : a[0:7] = 8'h2e;
            8'hbf : a[0:7] = 8'h20;
            8'hc0 : a[0:7] = 8'hec;
            8'hc1 : a[0:7] = 8'he2;
            8'hc2 : a[0:7] = 8'hf0;
            8'hc3 : a[0:7] = 8'hfe;
            8'hc4 : a[0:7] = 8'hd4;
            8'hc5 : a[0:7] = 8'hda;
            8'hc6 : a[0:7] = 8'hc8;
            8'hc7 : a[0:7] = 8'hc6;
            8'hc8 : a[0:7] = 8'h9c;
            8'hc9 : a[0:7] = 8'h92;
            8'hca : a[0:7] = 8'h80;
            8'hcb : a[0:7] = 8'h8e;
            8'hcc : a[0:7] = 8'ha4;
            8'hcd : a[0:7] = 8'haa;
            8'hce : a[0:7] = 8'hb8;
            8'hcf : a[0:7] = 8'hb6;
            8'hd0 : a[0:7] = 8'hc;
            8'hd1 : a[0:7] = 8'h2;
            8'hd2 : a[0:7] = 8'h10;
            8'hd3 : a[0:7] = 8'h1e;
            8'hd4 : a[0:7] = 8'h34;
            8'hd5 : a[0:7] = 8'h3a;
            8'hd6 : a[0:7] = 8'h28;
            8'hd7 : a[0:7] = 8'h26;
            8'hd8 : a[0:7] = 8'h7c;
            8'hd9 : a[0:7] = 8'h72;
            8'hda : a[0:7] = 8'h60;
            8'hdb : a[0:7] = 8'h6e;
            8'hdc : a[0:7] = 8'h44;
            8'hdd : a[0:7] = 8'h4a;
            8'hde : a[0:7] = 8'h58;
            8'hdf : a[0:7] = 8'h56;
            8'he0 : a[0:7] = 8'h37;
            8'he1 : a[0:7] = 8'h39;
            8'he2 : a[0:7] = 8'h2b;
            8'he3 : a[0:7] = 8'h25;
            8'he4 : a[0:7] = 8'hf;
            8'he5 : a[0:7] = 8'h1;
            8'he6 : a[0:7] = 8'h13;
            8'he7 : a[0:7] = 8'h1d;
            8'he8 : a[0:7] = 8'h47;
            8'he9 : a[0:7] = 8'h49;
            8'hea : a[0:7] = 8'h5b;
            8'heb : a[0:7] = 8'h55;
            8'hec : a[0:7] = 8'h7f;
            8'hed : a[0:7] = 8'h71;
            8'hee : a[0:7] = 8'h63;
            8'hef : a[0:7] = 8'h6d;
            8'hf0 : a[0:7] = 8'hd7;
            8'hf1 : a[0:7] = 8'hd9;
            8'hf2 : a[0:7] = 8'hcb;
            8'hf3 : a[0:7] = 8'hc5;
            8'hf4 : a[0:7] = 8'hef;
            8'hf5 : a[0:7] = 8'he1;
            8'hf6 : a[0:7] = 8'hf3;
            8'hf7 : a[0:7] = 8'hfd;
            8'hf8 : a[0:7] = 8'ha7;
            8'hf9 : a[0:7] = 8'ha9;
            8'hfa : a[0:7] = 8'hbb;
            8'hfb : a[0:7] = 8'hb5;
            8'hfc : a[0:7] = 8'h9f;
            8'hfd : a[0:7] = 8'h91;
            8'hfe : a[0:7] = 8'h83;
            8'hff : a[0:7] = 8'h8d;
        endcase
    end

    // Multiplication with 11
    always @(row[24:31]) begin
        case (row[24:31])
                        8'h0 : b[0:7] = 8'h0;
            8'h1 : b[0:7] = 8'hb;
            8'h2 : b[0:7] = 8'h16;
            8'h3 : b[0:7] = 8'h1d;
            8'h4 : b[0:7] = 8'h2c;
            8'h5 : b[0:7] = 8'h27;
            8'h6 : b[0:7] = 8'h3a;
            8'h7 : b[0:7] = 8'h31;
            8'h8 : b[0:7] = 8'h58;
            8'h9 : b[0:7] = 8'h53;
            8'ha : b[0:7] = 8'h4e;
            8'hb : b[0:7] = 8'h45;
            8'hc : b[0:7] = 8'h74;
            8'hd : b[0:7] = 8'h7f;
            8'he : b[0:7] = 8'h62;
            8'hf : b[0:7] = 8'h69;
            8'h10 : b[0:7] = 8'hb0;
            8'h11 : b[0:7] = 8'hbb;
            8'h12 : b[0:7] = 8'ha6;
            8'h13 : b[0:7] = 8'had;
            8'h14 : b[0:7] = 8'h9c;
            8'h15 : b[0:7] = 8'h97;
            8'h16 : b[0:7] = 8'h8a;
            8'h17 : b[0:7] = 8'h81;
            8'h18 : b[0:7] = 8'he8;
            8'h19 : b[0:7] = 8'he3;
            8'h1a : b[0:7] = 8'hfe;
            8'h1b : b[0:7] = 8'hf5;
            8'h1c : b[0:7] = 8'hc4;
            8'h1d : b[0:7] = 8'hcf;
            8'h1e : b[0:7] = 8'hd2;
            8'h1f : b[0:7] = 8'hd9;
            8'h20 : b[0:7] = 8'h7b;
            8'h21 : b[0:7] = 8'h70;
            8'h22 : b[0:7] = 8'h6d;
            8'h23 : b[0:7] = 8'h66;
            8'h24 : b[0:7] = 8'h57;
            8'h25 : b[0:7] = 8'h5c;
            8'h26 : b[0:7] = 8'h41;
            8'h27 : b[0:7] = 8'h4a;
            8'h28 : b[0:7] = 8'h23;
            8'h29 : b[0:7] = 8'h28;
            8'h2a : b[0:7] = 8'h35;
            8'h2b : b[0:7] = 8'h3e;
            8'h2c : b[0:7] = 8'hf;
            8'h2d : b[0:7] = 8'h4;
            8'h2e : b[0:7] = 8'h19;
            8'h2f : b[0:7] = 8'h12;
            8'h30 : b[0:7] = 8'hcb;
            8'h31 : b[0:7] = 8'hc0;
            8'h32 : b[0:7] = 8'hdd;
            8'h33 : b[0:7] = 8'hd6;
            8'h34 : b[0:7] = 8'he7;
            8'h35 : b[0:7] = 8'hec;
            8'h36 : b[0:7] = 8'hf1;
            8'h37 : b[0:7] = 8'hfa;
            8'h38 : b[0:7] = 8'h93;
            8'h39 : b[0:7] = 8'h98;
            8'h3a : b[0:7] = 8'h85;
            8'h3b : b[0:7] = 8'h8e;
            8'h3c : b[0:7] = 8'hbf;
            8'h3d : b[0:7] = 8'hb4;
            8'h3e : b[0:7] = 8'ha9;
            8'h3f : b[0:7] = 8'ha2;
            8'h40 : b[0:7] = 8'hf6;
            8'h41 : b[0:7] = 8'hfd;
            8'h42 : b[0:7] = 8'he0;
            8'h43 : b[0:7] = 8'heb;
            8'h44 : b[0:7] = 8'hda;
            8'h45 : b[0:7] = 8'hd1;
            8'h46 : b[0:7] = 8'hcc;
            8'h47 : b[0:7] = 8'hc7;
            8'h48 : b[0:7] = 8'hae;
            8'h49 : b[0:7] = 8'ha5;
            8'h4a : b[0:7] = 8'hb8;
            8'h4b : b[0:7] = 8'hb3;
            8'h4c : b[0:7] = 8'h82;
            8'h4d : b[0:7] = 8'h89;
            8'h4e : b[0:7] = 8'h94;
            8'h4f : b[0:7] = 8'h9f;
            8'h50 : b[0:7] = 8'h46;
            8'h51 : b[0:7] = 8'h4d;
            8'h52 : b[0:7] = 8'h50;
            8'h53 : b[0:7] = 8'h5b;
            8'h54 : b[0:7] = 8'h6a;
            8'h55 : b[0:7] = 8'h61;
            8'h56 : b[0:7] = 8'h7c;
            8'h57 : b[0:7] = 8'h77;
            8'h58 : b[0:7] = 8'h1e;
            8'h59 : b[0:7] = 8'h15;
            8'h5a : b[0:7] = 8'h8;
            8'h5b : b[0:7] = 8'h3;
            8'h5c : b[0:7] = 8'h32;
            8'h5d : b[0:7] = 8'h39;
            8'h5e : b[0:7] = 8'h24;
            8'h5f : b[0:7] = 8'h2f;
            8'h60 : b[0:7] = 8'h8d;
            8'h61 : b[0:7] = 8'h86;
            8'h62 : b[0:7] = 8'h9b;
            8'h63 : b[0:7] = 8'h90;
            8'h64 : b[0:7] = 8'ha1;
            8'h65 : b[0:7] = 8'haa;
            8'h66 : b[0:7] = 8'hb7;
            8'h67 : b[0:7] = 8'hbc;
            8'h68 : b[0:7] = 8'hd5;
            8'h69 : b[0:7] = 8'hde;
            8'h6a : b[0:7] = 8'hc3;
            8'h6b : b[0:7] = 8'hc8;
            8'h6c : b[0:7] = 8'hf9;
            8'h6d : b[0:7] = 8'hf2;
            8'h6e : b[0:7] = 8'hef;
            8'h6f : b[0:7] = 8'he4;
            8'h70 : b[0:7] = 8'h3d;
            8'h71 : b[0:7] = 8'h36;
            8'h72 : b[0:7] = 8'h2b;
            8'h73 : b[0:7] = 8'h20;
            8'h74 : b[0:7] = 8'h11;
            8'h75 : b[0:7] = 8'h1a;
            8'h76 : b[0:7] = 8'h7;
            8'h77 : b[0:7] = 8'hc;
            8'h78 : b[0:7] = 8'h65;
            8'h79 : b[0:7] = 8'h6e;
            8'h7a : b[0:7] = 8'h73;
            8'h7b : b[0:7] = 8'h78;
            8'h7c : b[0:7] = 8'h49;
            8'h7d : b[0:7] = 8'h42;
            8'h7e : b[0:7] = 8'h5f;
            8'h7f : b[0:7] = 8'h54;
            8'h80 : b[0:7] = 8'hf7;
            8'h81 : b[0:7] = 8'hfc;
            8'h82 : b[0:7] = 8'he1;
            8'h83 : b[0:7] = 8'hea;
            8'h84 : b[0:7] = 8'hdb;
            8'h85 : b[0:7] = 8'hd0;
            8'h86 : b[0:7] = 8'hcd;
            8'h87 : b[0:7] = 8'hc6;
            8'h88 : b[0:7] = 8'haf;
            8'h89 : b[0:7] = 8'ha4;
            8'h8a : b[0:7] = 8'hb9;
            8'h8b : b[0:7] = 8'hb2;
            8'h8c : b[0:7] = 8'h83;
            8'h8d : b[0:7] = 8'h88;
            8'h8e : b[0:7] = 8'h95;
            8'h8f : b[0:7] = 8'h9e;
            8'h90 : b[0:7] = 8'h47;
            8'h91 : b[0:7] = 8'h4c;
            8'h92 : b[0:7] = 8'h51;
            8'h93 : b[0:7] = 8'h5a;
            8'h94 : b[0:7] = 8'h6b;
            8'h95 : b[0:7] = 8'h60;
            8'h96 : b[0:7] = 8'h7d;
            8'h97 : b[0:7] = 8'h76;
            8'h98 : b[0:7] = 8'h1f;
            8'h99 : b[0:7] = 8'h14;
            8'h9a : b[0:7] = 8'h9;
            8'h9b : b[0:7] = 8'h2;
            8'h9c : b[0:7] = 8'h33;
            8'h9d : b[0:7] = 8'h38;
            8'h9e : b[0:7] = 8'h25;
            8'h9f : b[0:7] = 8'h2e;
            8'ha0 : b[0:7] = 8'h8c;
            8'ha1 : b[0:7] = 8'h87;
            8'ha2 : b[0:7] = 8'h9a;
            8'ha3 : b[0:7] = 8'h91;
            8'ha4 : b[0:7] = 8'ha0;
            8'ha5 : b[0:7] = 8'hab;
            8'ha6 : b[0:7] = 8'hb6;
            8'ha7 : b[0:7] = 8'hbd;
            8'ha8 : b[0:7] = 8'hd4;
            8'ha9 : b[0:7] = 8'hdf;
            8'haa : b[0:7] = 8'hc2;
            8'hab : b[0:7] = 8'hc9;
            8'hac : b[0:7] = 8'hf8;
            8'had : b[0:7] = 8'hf3;
            8'hae : b[0:7] = 8'hee;
            8'haf : b[0:7] = 8'he5;
            8'hb0 : b[0:7] = 8'h3c;
            8'hb1 : b[0:7] = 8'h37;
            8'hb2 : b[0:7] = 8'h2a;
            8'hb3 : b[0:7] = 8'h21;
            8'hb4 : b[0:7] = 8'h10;
            8'hb5 : b[0:7] = 8'h1b;
            8'hb6 : b[0:7] = 8'h6;
            8'hb7 : b[0:7] = 8'hd;
            8'hb8 : b[0:7] = 8'h64;
            8'hb9 : b[0:7] = 8'h6f;
            8'hba : b[0:7] = 8'h72;
            8'hbb : b[0:7] = 8'h79;
            8'hbc : b[0:7] = 8'h48;
            8'hbd : b[0:7] = 8'h43;
            8'hbe : b[0:7] = 8'h5e;
            8'hbf : b[0:7] = 8'h55;
            8'hc0 : b[0:7] = 8'h1;
            8'hc1 : b[0:7] = 8'ha;
            8'hc2 : b[0:7] = 8'h17;
            8'hc3 : b[0:7] = 8'h1c;
            8'hc4 : b[0:7] = 8'h2d;
            8'hc5 : b[0:7] = 8'h26;
            8'hc6 : b[0:7] = 8'h3b;
            8'hc7 : b[0:7] = 8'h30;
            8'hc8 : b[0:7] = 8'h59;
            8'hc9 : b[0:7] = 8'h52;
            8'hca : b[0:7] = 8'h4f;
            8'hcb : b[0:7] = 8'h44;
            8'hcc : b[0:7] = 8'h75;
            8'hcd : b[0:7] = 8'h7e;
            8'hce : b[0:7] = 8'h63;
            8'hcf : b[0:7] = 8'h68;
            8'hd0 : b[0:7] = 8'hb1;
            8'hd1 : b[0:7] = 8'hba;
            8'hd2 : b[0:7] = 8'ha7;
            8'hd3 : b[0:7] = 8'hac;
            8'hd4 : b[0:7] = 8'h9d;
            8'hd5 : b[0:7] = 8'h96;
            8'hd6 : b[0:7] = 8'h8b;
            8'hd7 : b[0:7] = 8'h80;
            8'hd8 : b[0:7] = 8'he9;
            8'hd9 : b[0:7] = 8'he2;
            8'hda : b[0:7] = 8'hff;
            8'hdb : b[0:7] = 8'hf4;
            8'hdc : b[0:7] = 8'hc5;
            8'hdd : b[0:7] = 8'hce;
            8'hde : b[0:7] = 8'hd3;
            8'hdf : b[0:7] = 8'hd8;
            8'he0 : b[0:7] = 8'h7a;
            8'he1 : b[0:7] = 8'h71;
            8'he2 : b[0:7] = 8'h6c;
            8'he3 : b[0:7] = 8'h67;
            8'he4 : b[0:7] = 8'h56;
            8'he5 : b[0:7] = 8'h5d;
            8'he6 : b[0:7] = 8'h40;
            8'he7 : b[0:7] = 8'h4b;
            8'he8 : b[0:7] = 8'h22;
            8'he9 : b[0:7] = 8'h29;
            8'hea : b[0:7] = 8'h34;
            8'heb : b[0:7] = 8'h3f;
            8'hec : b[0:7] = 8'he;
            8'hed : b[0:7] = 8'h5;
            8'hee : b[0:7] = 8'h18;
            8'hef : b[0:7] = 8'h13;
            8'hf0 : b[0:7] = 8'hca;
            8'hf1 : b[0:7] = 8'hc1;
            8'hf2 : b[0:7] = 8'hdc;
            8'hf3 : b[0:7] = 8'hd7;
            8'hf4 : b[0:7] = 8'he6;
            8'hf5 : b[0:7] = 8'hed;
            8'hf6 : b[0:7] = 8'hf0;
            8'hf7 : b[0:7] = 8'hfb;
            8'hf8 : b[0:7] = 8'h92;
            8'hf9 : b[0:7] = 8'h99;
            8'hfa : b[0:7] = 8'h84;
            8'hfb : b[0:7] = 8'h8f;
            8'hfc : b[0:7] = 8'hbe;
            8'hfd : b[0:7] = 8'hb5;
            8'hfe : b[0:7] = 8'ha8;
            8'hff : b[0:7] = 8'ha3;
        endcase
    end

    assign output_row = a ^ b ^ c ^ d;
    
endmodule


module MixColumn4RowInverse (
    input wire [0:31] row,
    output wire [0:7] output_row
);
    reg [0:7] a, b, c, d;

    // Multiplication with 11
    always @(row[0:7]) begin
        case (row[0:7])
                        8'h0 : b[0:7] = 8'h0;
            8'h1 : b[0:7] = 8'hb;
            8'h2 : b[0:7] = 8'h16;
            8'h3 : b[0:7] = 8'h1d;
            8'h4 : b[0:7] = 8'h2c;
            8'h5 : b[0:7] = 8'h27;
            8'h6 : b[0:7] = 8'h3a;
            8'h7 : b[0:7] = 8'h31;
            8'h8 : b[0:7] = 8'h58;
            8'h9 : b[0:7] = 8'h53;
            8'ha : b[0:7] = 8'h4e;
            8'hb : b[0:7] = 8'h45;
            8'hc : b[0:7] = 8'h74;
            8'hd : b[0:7] = 8'h7f;
            8'he : b[0:7] = 8'h62;
            8'hf : b[0:7] = 8'h69;
            8'h10 : b[0:7] = 8'hb0;
            8'h11 : b[0:7] = 8'hbb;
            8'h12 : b[0:7] = 8'ha6;
            8'h13 : b[0:7] = 8'had;
            8'h14 : b[0:7] = 8'h9c;
            8'h15 : b[0:7] = 8'h97;
            8'h16 : b[0:7] = 8'h8a;
            8'h17 : b[0:7] = 8'h81;
            8'h18 : b[0:7] = 8'he8;
            8'h19 : b[0:7] = 8'he3;
            8'h1a : b[0:7] = 8'hfe;
            8'h1b : b[0:7] = 8'hf5;
            8'h1c : b[0:7] = 8'hc4;
            8'h1d : b[0:7] = 8'hcf;
            8'h1e : b[0:7] = 8'hd2;
            8'h1f : b[0:7] = 8'hd9;
            8'h20 : b[0:7] = 8'h7b;
            8'h21 : b[0:7] = 8'h70;
            8'h22 : b[0:7] = 8'h6d;
            8'h23 : b[0:7] = 8'h66;
            8'h24 : b[0:7] = 8'h57;
            8'h25 : b[0:7] = 8'h5c;
            8'h26 : b[0:7] = 8'h41;
            8'h27 : b[0:7] = 8'h4a;
            8'h28 : b[0:7] = 8'h23;
            8'h29 : b[0:7] = 8'h28;
            8'h2a : b[0:7] = 8'h35;
            8'h2b : b[0:7] = 8'h3e;
            8'h2c : b[0:7] = 8'hf;
            8'h2d : b[0:7] = 8'h4;
            8'h2e : b[0:7] = 8'h19;
            8'h2f : b[0:7] = 8'h12;
            8'h30 : b[0:7] = 8'hcb;
            8'h31 : b[0:7] = 8'hc0;
            8'h32 : b[0:7] = 8'hdd;
            8'h33 : b[0:7] = 8'hd6;
            8'h34 : b[0:7] = 8'he7;
            8'h35 : b[0:7] = 8'hec;
            8'h36 : b[0:7] = 8'hf1;
            8'h37 : b[0:7] = 8'hfa;
            8'h38 : b[0:7] = 8'h93;
            8'h39 : b[0:7] = 8'h98;
            8'h3a : b[0:7] = 8'h85;
            8'h3b : b[0:7] = 8'h8e;
            8'h3c : b[0:7] = 8'hbf;
            8'h3d : b[0:7] = 8'hb4;
            8'h3e : b[0:7] = 8'ha9;
            8'h3f : b[0:7] = 8'ha2;
            8'h40 : b[0:7] = 8'hf6;
            8'h41 : b[0:7] = 8'hfd;
            8'h42 : b[0:7] = 8'he0;
            8'h43 : b[0:7] = 8'heb;
            8'h44 : b[0:7] = 8'hda;
            8'h45 : b[0:7] = 8'hd1;
            8'h46 : b[0:7] = 8'hcc;
            8'h47 : b[0:7] = 8'hc7;
            8'h48 : b[0:7] = 8'hae;
            8'h49 : b[0:7] = 8'ha5;
            8'h4a : b[0:7] = 8'hb8;
            8'h4b : b[0:7] = 8'hb3;
            8'h4c : b[0:7] = 8'h82;
            8'h4d : b[0:7] = 8'h89;
            8'h4e : b[0:7] = 8'h94;
            8'h4f : b[0:7] = 8'h9f;
            8'h50 : b[0:7] = 8'h46;
            8'h51 : b[0:7] = 8'h4d;
            8'h52 : b[0:7] = 8'h50;
            8'h53 : b[0:7] = 8'h5b;
            8'h54 : b[0:7] = 8'h6a;
            8'h55 : b[0:7] = 8'h61;
            8'h56 : b[0:7] = 8'h7c;
            8'h57 : b[0:7] = 8'h77;
            8'h58 : b[0:7] = 8'h1e;
            8'h59 : b[0:7] = 8'h15;
            8'h5a : b[0:7] = 8'h8;
            8'h5b : b[0:7] = 8'h3;
            8'h5c : b[0:7] = 8'h32;
            8'h5d : b[0:7] = 8'h39;
            8'h5e : b[0:7] = 8'h24;
            8'h5f : b[0:7] = 8'h2f;
            8'h60 : b[0:7] = 8'h8d;
            8'h61 : b[0:7] = 8'h86;
            8'h62 : b[0:7] = 8'h9b;
            8'h63 : b[0:7] = 8'h90;
            8'h64 : b[0:7] = 8'ha1;
            8'h65 : b[0:7] = 8'haa;
            8'h66 : b[0:7] = 8'hb7;
            8'h67 : b[0:7] = 8'hbc;
            8'h68 : b[0:7] = 8'hd5;
            8'h69 : b[0:7] = 8'hde;
            8'h6a : b[0:7] = 8'hc3;
            8'h6b : b[0:7] = 8'hc8;
            8'h6c : b[0:7] = 8'hf9;
            8'h6d : b[0:7] = 8'hf2;
            8'h6e : b[0:7] = 8'hef;
            8'h6f : b[0:7] = 8'he4;
            8'h70 : b[0:7] = 8'h3d;
            8'h71 : b[0:7] = 8'h36;
            8'h72 : b[0:7] = 8'h2b;
            8'h73 : b[0:7] = 8'h20;
            8'h74 : b[0:7] = 8'h11;
            8'h75 : b[0:7] = 8'h1a;
            8'h76 : b[0:7] = 8'h7;
            8'h77 : b[0:7] = 8'hc;
            8'h78 : b[0:7] = 8'h65;
            8'h79 : b[0:7] = 8'h6e;
            8'h7a : b[0:7] = 8'h73;
            8'h7b : b[0:7] = 8'h78;
            8'h7c : b[0:7] = 8'h49;
            8'h7d : b[0:7] = 8'h42;
            8'h7e : b[0:7] = 8'h5f;
            8'h7f : b[0:7] = 8'h54;
            8'h80 : b[0:7] = 8'hf7;
            8'h81 : b[0:7] = 8'hfc;
            8'h82 : b[0:7] = 8'he1;
            8'h83 : b[0:7] = 8'hea;
            8'h84 : b[0:7] = 8'hdb;
            8'h85 : b[0:7] = 8'hd0;
            8'h86 : b[0:7] = 8'hcd;
            8'h87 : b[0:7] = 8'hc6;
            8'h88 : b[0:7] = 8'haf;
            8'h89 : b[0:7] = 8'ha4;
            8'h8a : b[0:7] = 8'hb9;
            8'h8b : b[0:7] = 8'hb2;
            8'h8c : b[0:7] = 8'h83;
            8'h8d : b[0:7] = 8'h88;
            8'h8e : b[0:7] = 8'h95;
            8'h8f : b[0:7] = 8'h9e;
            8'h90 : b[0:7] = 8'h47;
            8'h91 : b[0:7] = 8'h4c;
            8'h92 : b[0:7] = 8'h51;
            8'h93 : b[0:7] = 8'h5a;
            8'h94 : b[0:7] = 8'h6b;
            8'h95 : b[0:7] = 8'h60;
            8'h96 : b[0:7] = 8'h7d;
            8'h97 : b[0:7] = 8'h76;
            8'h98 : b[0:7] = 8'h1f;
            8'h99 : b[0:7] = 8'h14;
            8'h9a : b[0:7] = 8'h9;
            8'h9b : b[0:7] = 8'h2;
            8'h9c : b[0:7] = 8'h33;
            8'h9d : b[0:7] = 8'h38;
            8'h9e : b[0:7] = 8'h25;
            8'h9f : b[0:7] = 8'h2e;
            8'ha0 : b[0:7] = 8'h8c;
            8'ha1 : b[0:7] = 8'h87;
            8'ha2 : b[0:7] = 8'h9a;
            8'ha3 : b[0:7] = 8'h91;
            8'ha4 : b[0:7] = 8'ha0;
            8'ha5 : b[0:7] = 8'hab;
            8'ha6 : b[0:7] = 8'hb6;
            8'ha7 : b[0:7] = 8'hbd;
            8'ha8 : b[0:7] = 8'hd4;
            8'ha9 : b[0:7] = 8'hdf;
            8'haa : b[0:7] = 8'hc2;
            8'hab : b[0:7] = 8'hc9;
            8'hac : b[0:7] = 8'hf8;
            8'had : b[0:7] = 8'hf3;
            8'hae : b[0:7] = 8'hee;
            8'haf : b[0:7] = 8'he5;
            8'hb0 : b[0:7] = 8'h3c;
            8'hb1 : b[0:7] = 8'h37;
            8'hb2 : b[0:7] = 8'h2a;
            8'hb3 : b[0:7] = 8'h21;
            8'hb4 : b[0:7] = 8'h10;
            8'hb5 : b[0:7] = 8'h1b;
            8'hb6 : b[0:7] = 8'h6;
            8'hb7 : b[0:7] = 8'hd;
            8'hb8 : b[0:7] = 8'h64;
            8'hb9 : b[0:7] = 8'h6f;
            8'hba : b[0:7] = 8'h72;
            8'hbb : b[0:7] = 8'h79;
            8'hbc : b[0:7] = 8'h48;
            8'hbd : b[0:7] = 8'h43;
            8'hbe : b[0:7] = 8'h5e;
            8'hbf : b[0:7] = 8'h55;
            8'hc0 : b[0:7] = 8'h1;
            8'hc1 : b[0:7] = 8'ha;
            8'hc2 : b[0:7] = 8'h17;
            8'hc3 : b[0:7] = 8'h1c;
            8'hc4 : b[0:7] = 8'h2d;
            8'hc5 : b[0:7] = 8'h26;
            8'hc6 : b[0:7] = 8'h3b;
            8'hc7 : b[0:7] = 8'h30;
            8'hc8 : b[0:7] = 8'h59;
            8'hc9 : b[0:7] = 8'h52;
            8'hca : b[0:7] = 8'h4f;
            8'hcb : b[0:7] = 8'h44;
            8'hcc : b[0:7] = 8'h75;
            8'hcd : b[0:7] = 8'h7e;
            8'hce : b[0:7] = 8'h63;
            8'hcf : b[0:7] = 8'h68;
            8'hd0 : b[0:7] = 8'hb1;
            8'hd1 : b[0:7] = 8'hba;
            8'hd2 : b[0:7] = 8'ha7;
            8'hd3 : b[0:7] = 8'hac;
            8'hd4 : b[0:7] = 8'h9d;
            8'hd5 : b[0:7] = 8'h96;
            8'hd6 : b[0:7] = 8'h8b;
            8'hd7 : b[0:7] = 8'h80;
            8'hd8 : b[0:7] = 8'he9;
            8'hd9 : b[0:7] = 8'he2;
            8'hda : b[0:7] = 8'hff;
            8'hdb : b[0:7] = 8'hf4;
            8'hdc : b[0:7] = 8'hc5;
            8'hdd : b[0:7] = 8'hce;
            8'hde : b[0:7] = 8'hd3;
            8'hdf : b[0:7] = 8'hd8;
            8'he0 : b[0:7] = 8'h7a;
            8'he1 : b[0:7] = 8'h71;
            8'he2 : b[0:7] = 8'h6c;
            8'he3 : b[0:7] = 8'h67;
            8'he4 : b[0:7] = 8'h56;
            8'he5 : b[0:7] = 8'h5d;
            8'he6 : b[0:7] = 8'h40;
            8'he7 : b[0:7] = 8'h4b;
            8'he8 : b[0:7] = 8'h22;
            8'he9 : b[0:7] = 8'h29;
            8'hea : b[0:7] = 8'h34;
            8'heb : b[0:7] = 8'h3f;
            8'hec : b[0:7] = 8'he;
            8'hed : b[0:7] = 8'h5;
            8'hee : b[0:7] = 8'h18;
            8'hef : b[0:7] = 8'h13;
            8'hf0 : b[0:7] = 8'hca;
            8'hf1 : b[0:7] = 8'hc1;
            8'hf2 : b[0:7] = 8'hdc;
            8'hf3 : b[0:7] = 8'hd7;
            8'hf4 : b[0:7] = 8'he6;
            8'hf5 : b[0:7] = 8'hed;
            8'hf6 : b[0:7] = 8'hf0;
            8'hf7 : b[0:7] = 8'hfb;
            8'hf8 : b[0:7] = 8'h92;
            8'hf9 : b[0:7] = 8'h99;
            8'hfa : b[0:7] = 8'h84;
            8'hfb : b[0:7] = 8'h8f;
            8'hfc : b[0:7] = 8'hbe;
            8'hfd : b[0:7] = 8'hb5;
            8'hfe : b[0:7] = 8'ha8;
            8'hff : b[0:7] = 8'ha3;
        endcase
    end

    // Multiplication with 13
    always @(row[8:15]) begin
        case (row[8:15])
            			8'h0 : c[0:7] = 8'h0;
			8'h1 : c[0:7] = 8'hd;
			8'h2 : c[0:7] = 8'h1a;
			8'h3 : c[0:7] = 8'h17;
			8'h4 : c[0:7] = 8'h34;
			8'h5 : c[0:7] = 8'h39;
			8'h6 : c[0:7] = 8'h2e;
			8'h7 : c[0:7] = 8'h23;
			8'h8 : c[0:7] = 8'h68;
			8'h9 : c[0:7] = 8'h65;
			8'ha : c[0:7] = 8'h72;
			8'hb : c[0:7] = 8'h7f;
			8'hc : c[0:7] = 8'h5c;
			8'hd : c[0:7] = 8'h51;
			8'he : c[0:7] = 8'h46;
			8'hf : c[0:7] = 8'h4b;
			8'h10 : c[0:7] = 8'hd0;
			8'h11 : c[0:7] = 8'hdd;
			8'h12 : c[0:7] = 8'hca;
			8'h13 : c[0:7] = 8'hc7;
			8'h14 : c[0:7] = 8'he4;
			8'h15 : c[0:7] = 8'he9;
			8'h16 : c[0:7] = 8'hfe;
			8'h17 : c[0:7] = 8'hf3;
			8'h18 : c[0:7] = 8'hb8;
			8'h19 : c[0:7] = 8'hb5;
			8'h1a : c[0:7] = 8'ha2;
			8'h1b : c[0:7] = 8'haf;
			8'h1c : c[0:7] = 8'h8c;
			8'h1d : c[0:7] = 8'h81;
			8'h1e : c[0:7] = 8'h96;
			8'h1f : c[0:7] = 8'h9b;
			8'h20 : c[0:7] = 8'hbb;
			8'h21 : c[0:7] = 8'hb6;
			8'h22 : c[0:7] = 8'ha1;
			8'h23 : c[0:7] = 8'hac;
			8'h24 : c[0:7] = 8'h8f;
			8'h25 : c[0:7] = 8'h82;
			8'h26 : c[0:7] = 8'h95;
			8'h27 : c[0:7] = 8'h98;
			8'h28 : c[0:7] = 8'hd3;
			8'h29 : c[0:7] = 8'hde;
			8'h2a : c[0:7] = 8'hc9;
			8'h2b : c[0:7] = 8'hc4;
			8'h2c : c[0:7] = 8'he7;
			8'h2d : c[0:7] = 8'hea;
			8'h2e : c[0:7] = 8'hfd;
			8'h2f : c[0:7] = 8'hf0;
			8'h30 : c[0:7] = 8'h6b;
			8'h31 : c[0:7] = 8'h66;
			8'h32 : c[0:7] = 8'h71;
			8'h33 : c[0:7] = 8'h7c;
			8'h34 : c[0:7] = 8'h5f;
			8'h35 : c[0:7] = 8'h52;
			8'h36 : c[0:7] = 8'h45;
			8'h37 : c[0:7] = 8'h48;
			8'h38 : c[0:7] = 8'h3;
			8'h39 : c[0:7] = 8'he;
			8'h3a : c[0:7] = 8'h19;
			8'h3b : c[0:7] = 8'h14;
			8'h3c : c[0:7] = 8'h37;
			8'h3d : c[0:7] = 8'h3a;
			8'h3e : c[0:7] = 8'h2d;
			8'h3f : c[0:7] = 8'h20;
			8'h40 : c[0:7] = 8'h6d;
			8'h41 : c[0:7] = 8'h60;
			8'h42 : c[0:7] = 8'h77;
			8'h43 : c[0:7] = 8'h7a;
			8'h44 : c[0:7] = 8'h59;
			8'h45 : c[0:7] = 8'h54;
			8'h46 : c[0:7] = 8'h43;
			8'h47 : c[0:7] = 8'h4e;
			8'h48 : c[0:7] = 8'h5;
			8'h49 : c[0:7] = 8'h8;
			8'h4a : c[0:7] = 8'h1f;
			8'h4b : c[0:7] = 8'h12;
			8'h4c : c[0:7] = 8'h31;
			8'h4d : c[0:7] = 8'h3c;
			8'h4e : c[0:7] = 8'h2b;
			8'h4f : c[0:7] = 8'h26;
			8'h50 : c[0:7] = 8'hbd;
			8'h51 : c[0:7] = 8'hb0;
			8'h52 : c[0:7] = 8'ha7;
			8'h53 : c[0:7] = 8'haa;
			8'h54 : c[0:7] = 8'h89;
			8'h55 : c[0:7] = 8'h84;
			8'h56 : c[0:7] = 8'h93;
			8'h57 : c[0:7] = 8'h9e;
			8'h58 : c[0:7] = 8'hd5;
			8'h59 : c[0:7] = 8'hd8;
			8'h5a : c[0:7] = 8'hcf;
			8'h5b : c[0:7] = 8'hc2;
			8'h5c : c[0:7] = 8'he1;
			8'h5d : c[0:7] = 8'hec;
			8'h5e : c[0:7] = 8'hfb;
			8'h5f : c[0:7] = 8'hf6;
			8'h60 : c[0:7] = 8'hd6;
			8'h61 : c[0:7] = 8'hdb;
			8'h62 : c[0:7] = 8'hcc;
			8'h63 : c[0:7] = 8'hc1;
			8'h64 : c[0:7] = 8'he2;
			8'h65 : c[0:7] = 8'hef;
			8'h66 : c[0:7] = 8'hf8;
			8'h67 : c[0:7] = 8'hf5;
			8'h68 : c[0:7] = 8'hbe;
			8'h69 : c[0:7] = 8'hb3;
			8'h6a : c[0:7] = 8'ha4;
			8'h6b : c[0:7] = 8'ha9;
			8'h6c : c[0:7] = 8'h8a;
			8'h6d : c[0:7] = 8'h87;
			8'h6e : c[0:7] = 8'h90;
			8'h6f : c[0:7] = 8'h9d;
			8'h70 : c[0:7] = 8'h6;
			8'h71 : c[0:7] = 8'hb;
			8'h72 : c[0:7] = 8'h1c;
			8'h73 : c[0:7] = 8'h11;
			8'h74 : c[0:7] = 8'h32;
			8'h75 : c[0:7] = 8'h3f;
			8'h76 : c[0:7] = 8'h28;
			8'h77 : c[0:7] = 8'h25;
			8'h78 : c[0:7] = 8'h6e;
			8'h79 : c[0:7] = 8'h63;
			8'h7a : c[0:7] = 8'h74;
			8'h7b : c[0:7] = 8'h79;
			8'h7c : c[0:7] = 8'h5a;
			8'h7d : c[0:7] = 8'h57;
			8'h7e : c[0:7] = 8'h40;
			8'h7f : c[0:7] = 8'h4d;
			8'h80 : c[0:7] = 8'hda;
			8'h81 : c[0:7] = 8'hd7;
			8'h82 : c[0:7] = 8'hc0;
			8'h83 : c[0:7] = 8'hcd;
			8'h84 : c[0:7] = 8'hee;
			8'h85 : c[0:7] = 8'he3;
			8'h86 : c[0:7] = 8'hf4;
			8'h87 : c[0:7] = 8'hf9;
			8'h88 : c[0:7] = 8'hb2;
			8'h89 : c[0:7] = 8'hbf;
			8'h8a : c[0:7] = 8'ha8;
			8'h8b : c[0:7] = 8'ha5;
			8'h8c : c[0:7] = 8'h86;
			8'h8d : c[0:7] = 8'h8b;
			8'h8e : c[0:7] = 8'h9c;
			8'h8f : c[0:7] = 8'h91;
			8'h90 : c[0:7] = 8'ha;
			8'h91 : c[0:7] = 8'h7;
			8'h92 : c[0:7] = 8'h10;
			8'h93 : c[0:7] = 8'h1d;
			8'h94 : c[0:7] = 8'h3e;
			8'h95 : c[0:7] = 8'h33;
			8'h96 : c[0:7] = 8'h24;
			8'h97 : c[0:7] = 8'h29;
			8'h98 : c[0:7] = 8'h62;
			8'h99 : c[0:7] = 8'h6f;
			8'h9a : c[0:7] = 8'h78;
			8'h9b : c[0:7] = 8'h75;
			8'h9c : c[0:7] = 8'h56;
			8'h9d : c[0:7] = 8'h5b;
			8'h9e : c[0:7] = 8'h4c;
			8'h9f : c[0:7] = 8'h41;
			8'ha0 : c[0:7] = 8'h61;
			8'ha1 : c[0:7] = 8'h6c;
			8'ha2 : c[0:7] = 8'h7b;
			8'ha3 : c[0:7] = 8'h76;
			8'ha4 : c[0:7] = 8'h55;
			8'ha5 : c[0:7] = 8'h58;
			8'ha6 : c[0:7] = 8'h4f;
			8'ha7 : c[0:7] = 8'h42;
			8'ha8 : c[0:7] = 8'h9;
			8'ha9 : c[0:7] = 8'h4;
			8'haa : c[0:7] = 8'h13;
			8'hab : c[0:7] = 8'h1e;
			8'hac : c[0:7] = 8'h3d;
			8'had : c[0:7] = 8'h30;
			8'hae : c[0:7] = 8'h27;
			8'haf : c[0:7] = 8'h2a;
			8'hb0 : c[0:7] = 8'hb1;
			8'hb1 : c[0:7] = 8'hbc;
			8'hb2 : c[0:7] = 8'hab;
			8'hb3 : c[0:7] = 8'ha6;
			8'hb4 : c[0:7] = 8'h85;
			8'hb5 : c[0:7] = 8'h88;
			8'hb6 : c[0:7] = 8'h9f;
			8'hb7 : c[0:7] = 8'h92;
			8'hb8 : c[0:7] = 8'hd9;
			8'hb9 : c[0:7] = 8'hd4;
			8'hba : c[0:7] = 8'hc3;
			8'hbb : c[0:7] = 8'hce;
			8'hbc : c[0:7] = 8'hed;
			8'hbd : c[0:7] = 8'he0;
			8'hbe : c[0:7] = 8'hf7;
			8'hbf : c[0:7] = 8'hfa;
			8'hc0 : c[0:7] = 8'hb7;
			8'hc1 : c[0:7] = 8'hba;
			8'hc2 : c[0:7] = 8'had;
			8'hc3 : c[0:7] = 8'ha0;
			8'hc4 : c[0:7] = 8'h83;
			8'hc5 : c[0:7] = 8'h8e;
			8'hc6 : c[0:7] = 8'h99;
			8'hc7 : c[0:7] = 8'h94;
			8'hc8 : c[0:7] = 8'hdf;
			8'hc9 : c[0:7] = 8'hd2;
			8'hca : c[0:7] = 8'hc5;
			8'hcb : c[0:7] = 8'hc8;
			8'hcc : c[0:7] = 8'heb;
			8'hcd : c[0:7] = 8'he6;
			8'hce : c[0:7] = 8'hf1;
			8'hcf : c[0:7] = 8'hfc;
			8'hd0 : c[0:7] = 8'h67;
			8'hd1 : c[0:7] = 8'h6a;
			8'hd2 : c[0:7] = 8'h7d;
			8'hd3 : c[0:7] = 8'h70;
			8'hd4 : c[0:7] = 8'h53;
			8'hd5 : c[0:7] = 8'h5e;
			8'hd6 : c[0:7] = 8'h49;
			8'hd7 : c[0:7] = 8'h44;
			8'hd8 : c[0:7] = 8'hf;
			8'hd9 : c[0:7] = 8'h2;
			8'hda : c[0:7] = 8'h15;
			8'hdb : c[0:7] = 8'h18;
			8'hdc : c[0:7] = 8'h3b;
			8'hdd : c[0:7] = 8'h36;
			8'hde : c[0:7] = 8'h21;
			8'hdf : c[0:7] = 8'h2c;
			8'he0 : c[0:7] = 8'hc;
			8'he1 : c[0:7] = 8'h1;
			8'he2 : c[0:7] = 8'h16;
			8'he3 : c[0:7] = 8'h1b;
			8'he4 : c[0:7] = 8'h38;
			8'he5 : c[0:7] = 8'h35;
			8'he6 : c[0:7] = 8'h22;
			8'he7 : c[0:7] = 8'h2f;
			8'he8 : c[0:7] = 8'h64;
			8'he9 : c[0:7] = 8'h69;
			8'hea : c[0:7] = 8'h7e;
			8'heb : c[0:7] = 8'h73;
			8'hec : c[0:7] = 8'h50;
			8'hed : c[0:7] = 8'h5d;
			8'hee : c[0:7] = 8'h4a;
			8'hef : c[0:7] = 8'h47;
			8'hf0 : c[0:7] = 8'hdc;
			8'hf1 : c[0:7] = 8'hd1;
			8'hf2 : c[0:7] = 8'hc6;
			8'hf3 : c[0:7] = 8'hcb;
			8'hf4 : c[0:7] = 8'he8;
			8'hf5 : c[0:7] = 8'he5;
			8'hf6 : c[0:7] = 8'hf2;
			8'hf7 : c[0:7] = 8'hff;
			8'hf8 : c[0:7] = 8'hb4;
			8'hf9 : c[0:7] = 8'hb9;
			8'hfa : c[0:7] = 8'hae;
			8'hfb : c[0:7] = 8'ha3;
			8'hfc : c[0:7] = 8'h80;
			8'hfd : c[0:7] = 8'h8d;
			8'hfe : c[0:7] = 8'h9a;
			8'hff : c[0:7] = 8'h97;
        endcase
    end

    // Multiplication with 9
    always @(row[16:23]) begin
        case (row[16:23])
			8'h0 : d[0:7] = 8'h0;
			8'h1 : d[0:7] = 8'h9;
			8'h2 : d[0:7] = 8'h12;
			8'h3 : d[0:7] = 8'h1b;
			8'h4 : d[0:7] = 8'h24;
			8'h5 : d[0:7] = 8'h2d;
			8'h6 : d[0:7] = 8'h36;
			8'h7 : d[0:7] = 8'h3f;
			8'h8 : d[0:7] = 8'h48;
			8'h9 : d[0:7] = 8'h41;
			8'ha : d[0:7] = 8'h5a;
			8'hb : d[0:7] = 8'h53;
			8'hc : d[0:7] = 8'h6c;
			8'hd : d[0:7] = 8'h65;
			8'he : d[0:7] = 8'h7e;
			8'hf : d[0:7] = 8'h77;
			8'h10 : d[0:7] = 8'h90;
			8'h11 : d[0:7] = 8'h99;
			8'h12 : d[0:7] = 8'h82;
			8'h13 : d[0:7] = 8'h8b;
			8'h14 : d[0:7] = 8'hb4;
			8'h15 : d[0:7] = 8'hbd;
			8'h16 : d[0:7] = 8'ha6;
			8'h17 : d[0:7] = 8'haf;
			8'h18 : d[0:7] = 8'hd8;
			8'h19 : d[0:7] = 8'hd1;
			8'h1a : d[0:7] = 8'hca;
			8'h1b : d[0:7] = 8'hc3;
			8'h1c : d[0:7] = 8'hfc;
			8'h1d : d[0:7] = 8'hf5;
			8'h1e : d[0:7] = 8'hee;
			8'h1f : d[0:7] = 8'he7;
			8'h20 : d[0:7] = 8'h3b;
			8'h21 : d[0:7] = 8'h32;
			8'h22 : d[0:7] = 8'h29;
			8'h23 : d[0:7] = 8'h20;
			8'h24 : d[0:7] = 8'h1f;
			8'h25 : d[0:7] = 8'h16;
			8'h26 : d[0:7] = 8'hd;
			8'h27 : d[0:7] = 8'h4;
			8'h28 : d[0:7] = 8'h73;
			8'h29 : d[0:7] = 8'h7a;
			8'h2a : d[0:7] = 8'h61;
			8'h2b : d[0:7] = 8'h68;
			8'h2c : d[0:7] = 8'h57;
			8'h2d : d[0:7] = 8'h5e;
			8'h2e : d[0:7] = 8'h45;
			8'h2f : d[0:7] = 8'h4c;
			8'h30 : d[0:7] = 8'hab;
			8'h31 : d[0:7] = 8'ha2;
			8'h32 : d[0:7] = 8'hb9;
			8'h33 : d[0:7] = 8'hb0;
			8'h34 : d[0:7] = 8'h8f;
			8'h35 : d[0:7] = 8'h86;
			8'h36 : d[0:7] = 8'h9d;
			8'h37 : d[0:7] = 8'h94;
			8'h38 : d[0:7] = 8'he3;
			8'h39 : d[0:7] = 8'hea;
			8'h3a : d[0:7] = 8'hf1;
			8'h3b : d[0:7] = 8'hf8;
			8'h3c : d[0:7] = 8'hc7;
			8'h3d : d[0:7] = 8'hce;
			8'h3e : d[0:7] = 8'hd5;
			8'h3f : d[0:7] = 8'hdc;
			8'h40 : d[0:7] = 8'h76;
			8'h41 : d[0:7] = 8'h7f;
			8'h42 : d[0:7] = 8'h64;
			8'h43 : d[0:7] = 8'h6d;
			8'h44 : d[0:7] = 8'h52;
			8'h45 : d[0:7] = 8'h5b;
			8'h46 : d[0:7] = 8'h40;
			8'h47 : d[0:7] = 8'h49;
			8'h48 : d[0:7] = 8'h3e;
			8'h49 : d[0:7] = 8'h37;
			8'h4a : d[0:7] = 8'h2c;
			8'h4b : d[0:7] = 8'h25;
			8'h4c : d[0:7] = 8'h1a;
			8'h4d : d[0:7] = 8'h13;
			8'h4e : d[0:7] = 8'h8;
			8'h4f : d[0:7] = 8'h1;
			8'h50 : d[0:7] = 8'he6;
			8'h51 : d[0:7] = 8'hef;
			8'h52 : d[0:7] = 8'hf4;
			8'h53 : d[0:7] = 8'hfd;
			8'h54 : d[0:7] = 8'hc2;
			8'h55 : d[0:7] = 8'hcb;
			8'h56 : d[0:7] = 8'hd0;
			8'h57 : d[0:7] = 8'hd9;
			8'h58 : d[0:7] = 8'hae;
			8'h59 : d[0:7] = 8'ha7;
			8'h5a : d[0:7] = 8'hbc;
			8'h5b : d[0:7] = 8'hb5;
			8'h5c : d[0:7] = 8'h8a;
			8'h5d : d[0:7] = 8'h83;
			8'h5e : d[0:7] = 8'h98;
			8'h5f : d[0:7] = 8'h91;
			8'h60 : d[0:7] = 8'h4d;
			8'h61 : d[0:7] = 8'h44;
			8'h62 : d[0:7] = 8'h5f;
			8'h63 : d[0:7] = 8'h56;
			8'h64 : d[0:7] = 8'h69;
			8'h65 : d[0:7] = 8'h60;
			8'h66 : d[0:7] = 8'h7b;
			8'h67 : d[0:7] = 8'h72;
			8'h68 : d[0:7] = 8'h5;
			8'h69 : d[0:7] = 8'hc;
			8'h6a : d[0:7] = 8'h17;
			8'h6b : d[0:7] = 8'h1e;
			8'h6c : d[0:7] = 8'h21;
			8'h6d : d[0:7] = 8'h28;
			8'h6e : d[0:7] = 8'h33;
			8'h6f : d[0:7] = 8'h3a;
			8'h70 : d[0:7] = 8'hdd;
			8'h71 : d[0:7] = 8'hd4;
			8'h72 : d[0:7] = 8'hcf;
			8'h73 : d[0:7] = 8'hc6;
			8'h74 : d[0:7] = 8'hf9;
			8'h75 : d[0:7] = 8'hf0;
			8'h76 : d[0:7] = 8'heb;
			8'h77 : d[0:7] = 8'he2;
			8'h78 : d[0:7] = 8'h95;
			8'h79 : d[0:7] = 8'h9c;
			8'h7a : d[0:7] = 8'h87;
			8'h7b : d[0:7] = 8'h8e;
			8'h7c : d[0:7] = 8'hb1;
			8'h7d : d[0:7] = 8'hb8;
			8'h7e : d[0:7] = 8'ha3;
			8'h7f : d[0:7] = 8'haa;
			8'h80 : d[0:7] = 8'hec;
			8'h81 : d[0:7] = 8'he5;
			8'h82 : d[0:7] = 8'hfe;
			8'h83 : d[0:7] = 8'hf7;
			8'h84 : d[0:7] = 8'hc8;
			8'h85 : d[0:7] = 8'hc1;
			8'h86 : d[0:7] = 8'hda;
			8'h87 : d[0:7] = 8'hd3;
			8'h88 : d[0:7] = 8'ha4;
			8'h89 : d[0:7] = 8'had;
			8'h8a : d[0:7] = 8'hb6;
			8'h8b : d[0:7] = 8'hbf;
			8'h8c : d[0:7] = 8'h80;
			8'h8d : d[0:7] = 8'h89;
			8'h8e : d[0:7] = 8'h92;
			8'h8f : d[0:7] = 8'h9b;
			8'h90 : d[0:7] = 8'h7c;
			8'h91 : d[0:7] = 8'h75;
			8'h92 : d[0:7] = 8'h6e;
			8'h93 : d[0:7] = 8'h67;
			8'h94 : d[0:7] = 8'h58;
			8'h95 : d[0:7] = 8'h51;
			8'h96 : d[0:7] = 8'h4a;
			8'h97 : d[0:7] = 8'h43;
			8'h98 : d[0:7] = 8'h34;
			8'h99 : d[0:7] = 8'h3d;
			8'h9a : d[0:7] = 8'h26;
			8'h9b : d[0:7] = 8'h2f;
			8'h9c : d[0:7] = 8'h10;
			8'h9d : d[0:7] = 8'h19;
			8'h9e : d[0:7] = 8'h2;
			8'h9f : d[0:7] = 8'hb;
			8'ha0 : d[0:7] = 8'hd7;
			8'ha1 : d[0:7] = 8'hde;
			8'ha2 : d[0:7] = 8'hc5;
			8'ha3 : d[0:7] = 8'hcc;
			8'ha4 : d[0:7] = 8'hf3;
			8'ha5 : d[0:7] = 8'hfa;
			8'ha6 : d[0:7] = 8'he1;
			8'ha7 : d[0:7] = 8'he8;
			8'ha8 : d[0:7] = 8'h9f;
			8'ha9 : d[0:7] = 8'h96;
			8'haa : d[0:7] = 8'h8d;
			8'hab : d[0:7] = 8'h84;
			8'hac : d[0:7] = 8'hbb;
			8'had : d[0:7] = 8'hb2;
			8'hae : d[0:7] = 8'ha9;
			8'haf : d[0:7] = 8'ha0;
			8'hb0 : d[0:7] = 8'h47;
			8'hb1 : d[0:7] = 8'h4e;
			8'hb2 : d[0:7] = 8'h55;
			8'hb3 : d[0:7] = 8'h5c;
			8'hb4 : d[0:7] = 8'h63;
			8'hb5 : d[0:7] = 8'h6a;
			8'hb6 : d[0:7] = 8'h71;
			8'hb7 : d[0:7] = 8'h78;
			8'hb8 : d[0:7] = 8'hf;
			8'hb9 : d[0:7] = 8'h6;
			8'hba : d[0:7] = 8'h1d;
			8'hbb : d[0:7] = 8'h14;
			8'hbc : d[0:7] = 8'h2b;
			8'hbd : d[0:7] = 8'h22;
			8'hbe : d[0:7] = 8'h39;
			8'hbf : d[0:7] = 8'h30;
			8'hc0 : d[0:7] = 8'h9a;
			8'hc1 : d[0:7] = 8'h93;
			8'hc2 : d[0:7] = 8'h88;
			8'hc3 : d[0:7] = 8'h81;
			8'hc4 : d[0:7] = 8'hbe;
			8'hc5 : d[0:7] = 8'hb7;
			8'hc6 : d[0:7] = 8'hac;
			8'hc7 : d[0:7] = 8'ha5;
			8'hc8 : d[0:7] = 8'hd2;
			8'hc9 : d[0:7] = 8'hdb;
			8'hca : d[0:7] = 8'hc0;
			8'hcb : d[0:7] = 8'hc9;
			8'hcc : d[0:7] = 8'hf6;
			8'hcd : d[0:7] = 8'hff;
			8'hce : d[0:7] = 8'he4;
			8'hcf : d[0:7] = 8'hed;
			8'hd0 : d[0:7] = 8'ha;
			8'hd1 : d[0:7] = 8'h3;
			8'hd2 : d[0:7] = 8'h18;
			8'hd3 : d[0:7] = 8'h11;
			8'hd4 : d[0:7] = 8'h2e;
			8'hd5 : d[0:7] = 8'h27;
			8'hd6 : d[0:7] = 8'h3c;
			8'hd7 : d[0:7] = 8'h35;
			8'hd8 : d[0:7] = 8'h42;
			8'hd9 : d[0:7] = 8'h4b;
			8'hda : d[0:7] = 8'h50;
			8'hdb : d[0:7] = 8'h59;
			8'hdc : d[0:7] = 8'h66;
			8'hdd : d[0:7] = 8'h6f;
			8'hde : d[0:7] = 8'h74;
			8'hdf : d[0:7] = 8'h7d;
			8'he0 : d[0:7] = 8'ha1;
			8'he1 : d[0:7] = 8'ha8;
			8'he2 : d[0:7] = 8'hb3;
			8'he3 : d[0:7] = 8'hba;
			8'he4 : d[0:7] = 8'h85;
			8'he5 : d[0:7] = 8'h8c;
			8'he6 : d[0:7] = 8'h97;
			8'he7 : d[0:7] = 8'h9e;
			8'he8 : d[0:7] = 8'he9;
			8'he9 : d[0:7] = 8'he0;
			8'hea : d[0:7] = 8'hfb;
			8'heb : d[0:7] = 8'hf2;
			8'hec : d[0:7] = 8'hcd;
			8'hed : d[0:7] = 8'hc4;
			8'hee : d[0:7] = 8'hdf;
			8'hef : d[0:7] = 8'hd6;
			8'hf0 : d[0:7] = 8'h31;
			8'hf1 : d[0:7] = 8'h38;
			8'hf2 : d[0:7] = 8'h23;
			8'hf3 : d[0:7] = 8'h2a;
			8'hf4 : d[0:7] = 8'h15;
			8'hf5 : d[0:7] = 8'h1c;
			8'hf6 : d[0:7] = 8'h7;
			8'hf7 : d[0:7] = 8'he;
			8'hf8 : d[0:7] = 8'h79;
			8'hf9 : d[0:7] = 8'h70;
			8'hfa : d[0:7] = 8'h6b;
			8'hfb : d[0:7] = 8'h62;
			8'hfc : d[0:7] = 8'h5d;
			8'hfd : d[0:7] = 8'h54;
			8'hfe : d[0:7] = 8'h4f;
			8'hff : d[0:7] = 8'h46;
        endcase
    end

    // Multiplication with 14
    always @(row[24:31]) begin
        case (row[24:31])
			            8'h0 : a[0:7] = 8'h0;
            8'h1 : a[0:7] = 8'he;
            8'h2 : a[0:7] = 8'h1c;
            8'h3 : a[0:7] = 8'h12;
            8'h4 : a[0:7] = 8'h38;
            8'h5 : a[0:7] = 8'h36;
            8'h6 : a[0:7] = 8'h24;
            8'h7 : a[0:7] = 8'h2a;
            8'h8 : a[0:7] = 8'h70;
            8'h9 : a[0:7] = 8'h7e;
            8'ha : a[0:7] = 8'h6c;
            8'hb : a[0:7] = 8'h62;
            8'hc : a[0:7] = 8'h48;
            8'hd : a[0:7] = 8'h46;
            8'he : a[0:7] = 8'h54;
            8'hf : a[0:7] = 8'h5a;
            8'h10 : a[0:7] = 8'he0;
            8'h11 : a[0:7] = 8'hee;
            8'h12 : a[0:7] = 8'hfc;
            8'h13 : a[0:7] = 8'hf2;
            8'h14 : a[0:7] = 8'hd8;
            8'h15 : a[0:7] = 8'hd6;
            8'h16 : a[0:7] = 8'hc4;
            8'h17 : a[0:7] = 8'hca;
            8'h18 : a[0:7] = 8'h90;
            8'h19 : a[0:7] = 8'h9e;
            8'h1a : a[0:7] = 8'h8c;
            8'h1b : a[0:7] = 8'h82;
            8'h1c : a[0:7] = 8'ha8;
            8'h1d : a[0:7] = 8'ha6;
            8'h1e : a[0:7] = 8'hb4;
            8'h1f : a[0:7] = 8'hba;
            8'h20 : a[0:7] = 8'hdb;
            8'h21 : a[0:7] = 8'hd5;
            8'h22 : a[0:7] = 8'hc7;
            8'h23 : a[0:7] = 8'hc9;
            8'h24 : a[0:7] = 8'he3;
            8'h25 : a[0:7] = 8'hed;
            8'h26 : a[0:7] = 8'hff;
            8'h27 : a[0:7] = 8'hf1;
            8'h28 : a[0:7] = 8'hab;
            8'h29 : a[0:7] = 8'ha5;
            8'h2a : a[0:7] = 8'hb7;
            8'h2b : a[0:7] = 8'hb9;
            8'h2c : a[0:7] = 8'h93;
            8'h2d : a[0:7] = 8'h9d;
            8'h2e : a[0:7] = 8'h8f;
            8'h2f : a[0:7] = 8'h81;
            8'h30 : a[0:7] = 8'h3b;
            8'h31 : a[0:7] = 8'h35;
            8'h32 : a[0:7] = 8'h27;
            8'h33 : a[0:7] = 8'h29;
            8'h34 : a[0:7] = 8'h3;
            8'h35 : a[0:7] = 8'hd;
            8'h36 : a[0:7] = 8'h1f;
            8'h37 : a[0:7] = 8'h11;
            8'h38 : a[0:7] = 8'h4b;
            8'h39 : a[0:7] = 8'h45;
            8'h3a : a[0:7] = 8'h57;
            8'h3b : a[0:7] = 8'h59;
            8'h3c : a[0:7] = 8'h73;
            8'h3d : a[0:7] = 8'h7d;
            8'h3e : a[0:7] = 8'h6f;
            8'h3f : a[0:7] = 8'h61;
            8'h40 : a[0:7] = 8'had;
            8'h41 : a[0:7] = 8'ha3;
            8'h42 : a[0:7] = 8'hb1;
            8'h43 : a[0:7] = 8'hbf;
            8'h44 : a[0:7] = 8'h95;
            8'h45 : a[0:7] = 8'h9b;
            8'h46 : a[0:7] = 8'h89;
            8'h47 : a[0:7] = 8'h87;
            8'h48 : a[0:7] = 8'hdd;
            8'h49 : a[0:7] = 8'hd3;
            8'h4a : a[0:7] = 8'hc1;
            8'h4b : a[0:7] = 8'hcf;
            8'h4c : a[0:7] = 8'he5;
            8'h4d : a[0:7] = 8'heb;
            8'h4e : a[0:7] = 8'hf9;
            8'h4f : a[0:7] = 8'hf7;
            8'h50 : a[0:7] = 8'h4d;
            8'h51 : a[0:7] = 8'h43;
            8'h52 : a[0:7] = 8'h51;
            8'h53 : a[0:7] = 8'h5f;
            8'h54 : a[0:7] = 8'h75;
            8'h55 : a[0:7] = 8'h7b;
            8'h56 : a[0:7] = 8'h69;
            8'h57 : a[0:7] = 8'h67;
            8'h58 : a[0:7] = 8'h3d;
            8'h59 : a[0:7] = 8'h33;
            8'h5a : a[0:7] = 8'h21;
            8'h5b : a[0:7] = 8'h2f;
            8'h5c : a[0:7] = 8'h5;
            8'h5d : a[0:7] = 8'hb;
            8'h5e : a[0:7] = 8'h19;
            8'h5f : a[0:7] = 8'h17;
            8'h60 : a[0:7] = 8'h76;
            8'h61 : a[0:7] = 8'h78;
            8'h62 : a[0:7] = 8'h6a;
            8'h63 : a[0:7] = 8'h64;
            8'h64 : a[0:7] = 8'h4e;
            8'h65 : a[0:7] = 8'h40;
            8'h66 : a[0:7] = 8'h52;
            8'h67 : a[0:7] = 8'h5c;
            8'h68 : a[0:7] = 8'h6;
            8'h69 : a[0:7] = 8'h8;
            8'h6a : a[0:7] = 8'h1a;
            8'h6b : a[0:7] = 8'h14;
            8'h6c : a[0:7] = 8'h3e;
            8'h6d : a[0:7] = 8'h30;
            8'h6e : a[0:7] = 8'h22;
            8'h6f : a[0:7] = 8'h2c;
            8'h70 : a[0:7] = 8'h96;
            8'h71 : a[0:7] = 8'h98;
            8'h72 : a[0:7] = 8'h8a;
            8'h73 : a[0:7] = 8'h84;
            8'h74 : a[0:7] = 8'hae;
            8'h75 : a[0:7] = 8'ha0;
            8'h76 : a[0:7] = 8'hb2;
            8'h77 : a[0:7] = 8'hbc;
            8'h78 : a[0:7] = 8'he6;
            8'h79 : a[0:7] = 8'he8;
            8'h7a : a[0:7] = 8'hfa;
            8'h7b : a[0:7] = 8'hf4;
            8'h7c : a[0:7] = 8'hde;
            8'h7d : a[0:7] = 8'hd0;
            8'h7e : a[0:7] = 8'hc2;
            8'h7f : a[0:7] = 8'hcc;
            8'h80 : a[0:7] = 8'h41;
            8'h81 : a[0:7] = 8'h4f;
            8'h82 : a[0:7] = 8'h5d;
            8'h83 : a[0:7] = 8'h53;
            8'h84 : a[0:7] = 8'h79;
            8'h85 : a[0:7] = 8'h77;
            8'h86 : a[0:7] = 8'h65;
            8'h87 : a[0:7] = 8'h6b;
            8'h88 : a[0:7] = 8'h31;
            8'h89 : a[0:7] = 8'h3f;
            8'h8a : a[0:7] = 8'h2d;
            8'h8b : a[0:7] = 8'h23;
            8'h8c : a[0:7] = 8'h9;
            8'h8d : a[0:7] = 8'h7;
            8'h8e : a[0:7] = 8'h15;
            8'h8f : a[0:7] = 8'h1b;
            8'h90 : a[0:7] = 8'ha1;
            8'h91 : a[0:7] = 8'haf;
            8'h92 : a[0:7] = 8'hbd;
            8'h93 : a[0:7] = 8'hb3;
            8'h94 : a[0:7] = 8'h99;
            8'h95 : a[0:7] = 8'h97;
            8'h96 : a[0:7] = 8'h85;
            8'h97 : a[0:7] = 8'h8b;
            8'h98 : a[0:7] = 8'hd1;
            8'h99 : a[0:7] = 8'hdf;
            8'h9a : a[0:7] = 8'hcd;
            8'h9b : a[0:7] = 8'hc3;
            8'h9c : a[0:7] = 8'he9;
            8'h9d : a[0:7] = 8'he7;
            8'h9e : a[0:7] = 8'hf5;
            8'h9f : a[0:7] = 8'hfb;
            8'ha0 : a[0:7] = 8'h9a;
            8'ha1 : a[0:7] = 8'h94;
            8'ha2 : a[0:7] = 8'h86;
            8'ha3 : a[0:7] = 8'h88;
            8'ha4 : a[0:7] = 8'ha2;
            8'ha5 : a[0:7] = 8'hac;
            8'ha6 : a[0:7] = 8'hbe;
            8'ha7 : a[0:7] = 8'hb0;
            8'ha8 : a[0:7] = 8'hea;
            8'ha9 : a[0:7] = 8'he4;
            8'haa : a[0:7] = 8'hf6;
            8'hab : a[0:7] = 8'hf8;
            8'hac : a[0:7] = 8'hd2;
            8'had : a[0:7] = 8'hdc;
            8'hae : a[0:7] = 8'hce;
            8'haf : a[0:7] = 8'hc0;
            8'hb0 : a[0:7] = 8'h7a;
            8'hb1 : a[0:7] = 8'h74;
            8'hb2 : a[0:7] = 8'h66;
            8'hb3 : a[0:7] = 8'h68;
            8'hb4 : a[0:7] = 8'h42;
            8'hb5 : a[0:7] = 8'h4c;
            8'hb6 : a[0:7] = 8'h5e;
            8'hb7 : a[0:7] = 8'h50;
            8'hb8 : a[0:7] = 8'ha;
            8'hb9 : a[0:7] = 8'h4;
            8'hba : a[0:7] = 8'h16;
            8'hbb : a[0:7] = 8'h18;
            8'hbc : a[0:7] = 8'h32;
            8'hbd : a[0:7] = 8'h3c;
            8'hbe : a[0:7] = 8'h2e;
            8'hbf : a[0:7] = 8'h20;
            8'hc0 : a[0:7] = 8'hec;
            8'hc1 : a[0:7] = 8'he2;
            8'hc2 : a[0:7] = 8'hf0;
            8'hc3 : a[0:7] = 8'hfe;
            8'hc4 : a[0:7] = 8'hd4;
            8'hc5 : a[0:7] = 8'hda;
            8'hc6 : a[0:7] = 8'hc8;
            8'hc7 : a[0:7] = 8'hc6;
            8'hc8 : a[0:7] = 8'h9c;
            8'hc9 : a[0:7] = 8'h92;
            8'hca : a[0:7] = 8'h80;
            8'hcb : a[0:7] = 8'h8e;
            8'hcc : a[0:7] = 8'ha4;
            8'hcd : a[0:7] = 8'haa;
            8'hce : a[0:7] = 8'hb8;
            8'hcf : a[0:7] = 8'hb6;
            8'hd0 : a[0:7] = 8'hc;
            8'hd1 : a[0:7] = 8'h2;
            8'hd2 : a[0:7] = 8'h10;
            8'hd3 : a[0:7] = 8'h1e;
            8'hd4 : a[0:7] = 8'h34;
            8'hd5 : a[0:7] = 8'h3a;
            8'hd6 : a[0:7] = 8'h28;
            8'hd7 : a[0:7] = 8'h26;
            8'hd8 : a[0:7] = 8'h7c;
            8'hd9 : a[0:7] = 8'h72;
            8'hda : a[0:7] = 8'h60;
            8'hdb : a[0:7] = 8'h6e;
            8'hdc : a[0:7] = 8'h44;
            8'hdd : a[0:7] = 8'h4a;
            8'hde : a[0:7] = 8'h58;
            8'hdf : a[0:7] = 8'h56;
            8'he0 : a[0:7] = 8'h37;
            8'he1 : a[0:7] = 8'h39;
            8'he2 : a[0:7] = 8'h2b;
            8'he3 : a[0:7] = 8'h25;
            8'he4 : a[0:7] = 8'hf;
            8'he5 : a[0:7] = 8'h1;
            8'he6 : a[0:7] = 8'h13;
            8'he7 : a[0:7] = 8'h1d;
            8'he8 : a[0:7] = 8'h47;
            8'he9 : a[0:7] = 8'h49;
            8'hea : a[0:7] = 8'h5b;
            8'heb : a[0:7] = 8'h55;
            8'hec : a[0:7] = 8'h7f;
            8'hed : a[0:7] = 8'h71;
            8'hee : a[0:7] = 8'h63;
            8'hef : a[0:7] = 8'h6d;
            8'hf0 : a[0:7] = 8'hd7;
            8'hf1 : a[0:7] = 8'hd9;
            8'hf2 : a[0:7] = 8'hcb;
            8'hf3 : a[0:7] = 8'hc5;
            8'hf4 : a[0:7] = 8'hef;
            8'hf5 : a[0:7] = 8'he1;
            8'hf6 : a[0:7] = 8'hf3;
            8'hf7 : a[0:7] = 8'hfd;
            8'hf8 : a[0:7] = 8'ha7;
            8'hf9 : a[0:7] = 8'ha9;
            8'hfa : a[0:7] = 8'hbb;
            8'hfb : a[0:7] = 8'hb5;
            8'hfc : a[0:7] = 8'h9f;
            8'hfd : a[0:7] = 8'h91;
            8'hfe : a[0:7] = 8'h83;
            8'hff : a[0:7] = 8'h8d;			
        endcase
    end

    assign output_row = a ^ b ^ c ^ d;
    
endmodule


module MixColumnInverse (
    input wire [0:31] row,
    output wire [0:31] output_row
);
    wire [0:7] a, b, c, d;

    MixColumn1RowInverse MixColumn1RowInverseModule(row[0:31], a[0:7]);
    MixColumn2RowInverse MixColumn2RowInverseModule(row[0:31], b[0:7]);
    MixColumn3RowInverse MixColumn3RowInverseModule(row[0:31], c[0:7]);
    MixColumn4RowInverse MixColumn4RowInverseModule(row[0:31], d[0:7]);

    assign output_row[0:7] = a[0:7];
    assign output_row[8:15] = b[0:7];
    assign output_row[16:23] = c[0:7];
    assign output_row[24:31] = d[0:7];
    

    
endmodule