module subWord (
    input wire [0:7] w_in,
    output reg [0:7] w_out
);

    always @(w_in[0:7]) begin
        case(w_in[0:7])
            32'h0 : w_out = 32'h63;
            32'h1 : w_out = 32'h7C;
            32'h2 : w_out = 32'h77;
            32'h3 : w_out = 32'h7B;
            32'h4 : w_out = 32'hF2;
            32'h5 : w_out = 32'h6B;
            32'h6 : w_out = 32'h6F;
            32'h7 : w_out = 32'hC5;
            32'h8 : w_out = 32'h30;
            32'h9 : w_out = 32'h1;
            32'hA : w_out = 32'h67;
            32'hB : w_out = 32'h2B;
            32'hC : w_out = 32'hFE;
            32'hD : w_out = 32'hD7;
            32'hE : w_out = 32'hAB;
            32'hF : w_out = 32'h76;
            32'h10 : w_out = 32'hCA;
            32'h11 : w_out = 32'h82;
            32'h12 : w_out = 32'hC9;
            32'h13 : w_out = 32'h7D;
            32'h14 : w_out = 32'hFA;
            32'h15 : w_out = 32'h59;
            32'h16 : w_out = 32'h47;
            32'h17 : w_out = 32'hF0;
            32'h18 : w_out = 32'hAD;
            32'h19 : w_out = 32'hD4;
            32'h1A : w_out = 32'hA2;
            32'h1B : w_out = 32'hAF;
            32'h1C : w_out = 32'h9C;
            32'h1D : w_out = 32'hA4;
            32'h1E : w_out = 32'h72;
            32'h1F : w_out = 32'hC0;
            32'h20 : w_out = 32'hB7;
            32'h21 : w_out = 32'hFD;
            32'h22 : w_out = 32'h93;
            32'h23 : w_out = 32'h26;
            32'h24 : w_out = 32'h36;
            32'h25 : w_out = 32'h3F;
            32'h26 : w_out = 32'hF7;
            32'h27 : w_out = 32'hCC;
            32'h28 : w_out = 32'h34;
            32'h29 : w_out = 32'hA5;
            32'h2A : w_out = 32'hE5;
            32'h2B : w_out = 32'hF1;
            32'h2C : w_out = 32'h71;
            32'h2D : w_out = 32'hD8;
            32'h2E : w_out = 32'h31;
            32'h2F : w_out = 32'h15;
            32'h30 : w_out = 32'h4;
            32'h31 : w_out = 32'hC7;
            32'h32 : w_out = 32'h23;
            32'h33 : w_out = 32'hC3;
            32'h34 : w_out = 32'h18;
            32'h35 : w_out = 32'h96;
            32'h36 : w_out = 32'h5;
            32'h37 : w_out = 32'h9A;
            32'h38 : w_out = 32'h7;
            32'h39 : w_out = 32'h12;
            32'h3A : w_out = 32'h80;
            32'h3B : w_out = 32'hE2;
            32'h3C : w_out = 32'hEB;
            32'h3D : w_out = 32'h27;
            32'h3E : w_out = 32'hB2;
            32'h3F : w_out = 32'h75;
            32'h40 : w_out = 32'h9;
            32'h41 : w_out = 32'h83;
            32'h42 : w_out = 32'h2C;
            32'h43 : w_out = 32'h1A;
            32'h44 : w_out = 32'h1B;
            32'h45 : w_out = 32'h6E;
            32'h46 : w_out = 32'h5A;
            32'h47 : w_out = 32'hA0;
            32'h48 : w_out = 32'h52;
            32'h49 : w_out = 32'h3B;
            32'h4A : w_out = 32'hD6;
            32'h4B : w_out = 32'hB3;
            32'h4C : w_out = 32'h29;
            32'h4D : w_out = 32'hE3;
            32'h4E : w_out = 32'h2F;
            32'h4F : w_out = 32'h84;
            32'h50 : w_out = 32'h53;
            32'h51 : w_out = 32'hD1;
            32'h52 : w_out = 32'h0;
            32'h53 : w_out = 32'hED;
            32'h54 : w_out = 32'h20;
            32'h55 : w_out = 32'hFC;
            32'h56 : w_out = 32'hB1;
            32'h57 : w_out = 32'h5B;
            32'h58 : w_out = 32'h6A;
            32'h59 : w_out = 32'hCB;
            32'h5A : w_out = 32'hBE;
            32'h5B : w_out = 32'h39;
            32'h5C : w_out = 32'h4A;
            32'h5D : w_out = 32'h4C;
            32'h5E : w_out = 32'h58;
            32'h5F : w_out = 32'hCF;
            32'h60 : w_out = 32'hD0;
            32'h61 : w_out = 32'hEF;
            32'h62 : w_out = 32'hAA;
            32'h63 : w_out = 32'hFB;
            32'h64 : w_out = 32'h43;
            32'h65 : w_out = 32'h4D;
            32'h66 : w_out = 32'h33;
            32'h67 : w_out = 32'h85;
            32'h68 : w_out = 32'h45;
            32'h69 : w_out = 32'hF9;
            32'h6A : w_out = 32'h2;
            32'h6B : w_out = 32'h7F;
            32'h6C : w_out = 32'h50;
            32'h6D : w_out = 32'h3C;
            32'h6E : w_out = 32'h9F;
            32'h6F : w_out = 32'hA8;
            32'h70 : w_out = 32'h51;
            32'h71 : w_out = 32'hA3;
            32'h72 : w_out = 32'h40;
            32'h73 : w_out = 32'h8F;
            32'h74 : w_out = 32'h92;
            32'h75 : w_out = 32'h9D;
            32'h76 : w_out = 32'h38;
            32'h77 : w_out = 32'hF5;
            32'h78 : w_out = 32'hBC;
            32'h79 : w_out = 32'hB6;
            32'h7A : w_out = 32'hDA;
            32'h7B : w_out = 32'h21;
            32'h7C : w_out = 32'h10;
            32'h7D : w_out = 32'hFF;
            32'h7E : w_out = 32'hF3;
            32'h7F : w_out = 32'hD2;
            32'h80 : w_out = 32'hCD;
            32'h81 : w_out = 32'hC;
            32'h82 : w_out = 32'h13;
            32'h83 : w_out = 32'hEC;
            32'h84 : w_out = 32'h5F;
            32'h85 : w_out = 32'h97;
            32'h86 : w_out = 32'h44;
            32'h87 : w_out = 32'h17;
            32'h88 : w_out = 32'hC4;
            32'h89 : w_out = 32'hA7;
            32'h8A : w_out = 32'h7E;
            32'h8B : w_out = 32'h3D;
            32'h8C : w_out = 32'h64;
            32'h8D : w_out = 32'h5D;
            32'h8E : w_out = 32'h19;
            32'h8F : w_out = 32'h73;
            32'h90 : w_out = 32'h60;
            32'h91 : w_out = 32'h81;
            32'h92 : w_out = 32'h4F;
            32'h93 : w_out = 32'hDC;
            32'h94 : w_out = 32'h22;
            32'h95 : w_out = 32'h2A;
            32'h96 : w_out = 32'h90;
            32'h97 : w_out = 32'h88;
            32'h98 : w_out = 32'h46;
            32'h99 : w_out = 32'hEE;
            32'h9A : w_out = 32'hB8;
            32'h9B : w_out = 32'h14;
            32'h9C : w_out = 32'hDE;
            32'h9D : w_out = 32'h5E;
            32'h9E : w_out = 32'hB;
            32'h9F : w_out = 32'hDB;
            32'hA0 : w_out = 32'hE0;
            32'hA1 : w_out = 32'h32;
            32'hA2 : w_out = 32'h3A;
            32'hA3 : w_out = 32'hA;
            32'hA4 : w_out = 32'h49;
            32'hA5 : w_out = 32'h6;
            32'hA6 : w_out = 32'h24;
            32'hA7 : w_out = 32'h5C;
            32'hA8 : w_out = 32'hC2;
            32'hA9 : w_out = 32'hD3;
            32'hAA : w_out = 32'hAC;
            32'hAB : w_out = 32'h62;
            32'hAC : w_out = 32'h91;
            32'hAD : w_out = 32'h95;
            32'hAE : w_out = 32'hE4;
            32'hAF : w_out = 32'h79;
            32'hB0 : w_out = 32'hE7;
            32'hB1 : w_out = 32'hC8;
            32'hB2 : w_out = 32'h37;
            32'hB3 : w_out = 32'h6D;
            32'hB4 : w_out = 32'h8D;
            32'hB5 : w_out = 32'hD5;
            32'hB6 : w_out = 32'h4E;
            32'hB7 : w_out = 32'hA9;
            32'hB8 : w_out = 32'h6C;
            32'hB9 : w_out = 32'h56;
            32'hBA : w_out = 32'hF4;
            32'hBB : w_out = 32'hEA;
            32'hBC : w_out = 32'h65;
            32'hBD : w_out = 32'h7A;
            32'hBE : w_out = 32'hAE;
            32'hBF : w_out = 32'h8;
            32'hC0 : w_out = 32'hBA;
            32'hC1 : w_out = 32'h78;
            32'hC2 : w_out = 32'h25;
            32'hC3 : w_out = 32'h2E;
            32'hC4 : w_out = 32'h1C;
            32'hC5 : w_out = 32'hA6;
            32'hC6 : w_out = 32'hB4;
            32'hC7 : w_out = 32'hC6;
            32'hC8 : w_out = 32'hE8;
            32'hC9 : w_out = 32'hDD;
            32'hCA : w_out = 32'h74;
            32'hCB : w_out = 32'h1F;
            32'hCC : w_out = 32'h4B;
            32'hCD : w_out = 32'hBD;
            32'hCE : w_out = 32'h8B;
            32'hCF : w_out = 32'h8A;
            32'hD0 : w_out = 32'h70;
            32'hD1 : w_out = 32'h3E;
            32'hD2 : w_out = 32'hB5;
            32'hD3 : w_out = 32'h66;
            32'hD4 : w_out = 32'h48;
            32'hD5 : w_out = 32'h3;
            32'hD6 : w_out = 32'hF6;
            32'hD7 : w_out = 32'hE;
            32'hD8 : w_out = 32'h61;
            32'hD9 : w_out = 32'h35;
            32'hDA : w_out = 32'h57;
            32'hDB : w_out = 32'hB9;
            32'hDC : w_out = 32'h86;
            32'hDD : w_out = 32'hC1;
            32'hDE : w_out = 32'h1D;
            32'hDF : w_out = 32'h9E;
            32'hE0 : w_out = 32'hE1;
            32'hE1 : w_out = 32'hF8;
            32'hE2 : w_out = 32'h98;
            32'hE3 : w_out = 32'h11;
            32'hE4 : w_out = 32'h69;
            32'hE5 : w_out = 32'hD9;
            32'hE6 : w_out = 32'h8E;
            32'hE7 : w_out = 32'h94;
            32'hE8 : w_out = 32'h9B;
            32'hE9 : w_out = 32'h1E;
            32'hEA : w_out = 32'h87;
            32'hEB : w_out = 32'hE9;
            32'hEC : w_out = 32'hCE;
            32'hED : w_out = 32'h55;
            32'hEE : w_out = 32'h28;
            32'hEF : w_out = 32'hDF;
            32'hF0 : w_out = 32'h8C;
            32'hF1 : w_out = 32'hA1;
            32'hF2 : w_out = 32'h89;
            32'hF3 : w_out = 32'hD;
            32'hF4 : w_out = 32'hBF;
            32'hF5 : w_out = 32'hE6;
            32'hF6 : w_out = 32'h42;
            32'hF7 : w_out = 32'h68;
            32'hF8 : w_out = 32'h41;
            32'hF9 : w_out = 32'h99;
            32'hFA : w_out = 32'h2D;
            32'hFB : w_out = 32'hF;
            32'hFC : w_out = 32'hB0;
            32'hFD : w_out = 32'h54;
            32'hFE : w_out = 32'hBB;
            32'hFF : w_out = 32'h16;
        endcase
    end
    
endmodule