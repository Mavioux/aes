module MixColumn1Row (
    input wire [0:31] row,
    output wire [0:7] output_row
);
    reg [0:7] a, b, c, d;

    // Multiplication with 2
    always @(row[0:7]) begin
        case (row[0:7])
            8'h0 : a[0:7] = 8'h0;
            8'h1 : a[0:7] = 8'h2;
            8'h2 : a[0:7] = 8'h4;
            8'h3 : a[0:7] = 8'h6;
            8'h4 : a[0:7] = 8'h8;
            8'h5 : a[0:7] = 8'hA;
            8'h6 : a[0:7] = 8'hC;
            8'h7 : a[0:7] = 8'hE;
            8'h8 : a[0:7] = 8'h10;
            8'h9 : a[0:7] = 8'h12;
            8'hA : a[0:7] = 8'h14;
            8'hB : a[0:7] = 8'h16;
            8'hC : a[0:7] = 8'h18;
            8'hD : a[0:7] = 8'h1A;
            8'hE : a[0:7] = 8'h1C;
            8'hF : a[0:7] = 8'h1E;
            8'h10 : a[0:7] = 8'h20;
            8'h11 : a[0:7] = 8'h22;
            8'h12 : a[0:7] = 8'h24;
            8'h13 : a[0:7] = 8'h26;
            8'h14 : a[0:7] = 8'h28;
            8'h15 : a[0:7] = 8'h2A;
            8'h16 : a[0:7] = 8'h2C;
            8'h17 : a[0:7] = 8'h2E;
            8'h18 : a[0:7] = 8'h30;
            8'h19 : a[0:7] = 8'h32;
            8'h1A : a[0:7] = 8'h34;
            8'h1B : a[0:7] = 8'h36;
            8'h1C : a[0:7] = 8'h38;
            8'h1D : a[0:7] = 8'h3A;
            8'h1E : a[0:7] = 8'h3C;
            8'h1F : a[0:7] = 8'h3E;
            8'h20 : a[0:7] = 8'h40;
            8'h21 : a[0:7] = 8'h42;
            8'h22 : a[0:7] = 8'h44;
            8'h23 : a[0:7] = 8'h46;
            8'h24 : a[0:7] = 8'h48;
            8'h25 : a[0:7] = 8'h4A;
            8'h26 : a[0:7] = 8'h4C;
            8'h27 : a[0:7] = 8'h4E;
            8'h28 : a[0:7] = 8'h50;
            8'h29 : a[0:7] = 8'h52;
            8'h2A : a[0:7] = 8'h54;
            8'h2B : a[0:7] = 8'h56;
            8'h2C : a[0:7] = 8'h58;
            8'h2D : a[0:7] = 8'h5A;
            8'h2E : a[0:7] = 8'h5C;
            8'h2F : a[0:7] = 8'h5E;
            8'h30 : a[0:7] = 8'h60;
            8'h31 : a[0:7] = 8'h62;
            8'h32 : a[0:7] = 8'h64;
            8'h33 : a[0:7] = 8'h66;
            8'h34 : a[0:7] = 8'h68;
            8'h35 : a[0:7] = 8'h6A;
            8'h36 : a[0:7] = 8'h6C;
            8'h37 : a[0:7] = 8'h6E;
            8'h38 : a[0:7] = 8'h70;
            8'h39 : a[0:7] = 8'h72;
            8'h3A : a[0:7] = 8'h74;
            8'h3B : a[0:7] = 8'h76;
            8'h3C : a[0:7] = 8'h78;
            8'h3D : a[0:7] = 8'h7A;
            8'h3E : a[0:7] = 8'h7C;
            8'h3F : a[0:7] = 8'h7E;
            8'h40 : a[0:7] = 8'h80;
            8'h41 : a[0:7] = 8'h82;
            8'h42 : a[0:7] = 8'h84;
            8'h43 : a[0:7] = 8'h86;
            8'h44 : a[0:7] = 8'h88;
            8'h45 : a[0:7] = 8'h8A;
            8'h46 : a[0:7] = 8'h8C;
            8'h47 : a[0:7] = 8'h8E;
            8'h48 : a[0:7] = 8'h90;
            8'h49 : a[0:7] = 8'h92;
            8'h4A : a[0:7] = 8'h94;
            8'h4B : a[0:7] = 8'h96;
            8'h4C : a[0:7] = 8'h98;
            8'h4D : a[0:7] = 8'h9A;
            8'h4E : a[0:7] = 8'h9C;
            8'h4F : a[0:7] = 8'h9E;
            8'h50 : a[0:7] = 8'hA0;
            8'h51 : a[0:7] = 8'hA2;
            8'h52 : a[0:7] = 8'hA4;
            8'h53 : a[0:7] = 8'hA6;
            8'h54 : a[0:7] = 8'hA8;
            8'h55 : a[0:7] = 8'hAA;
            8'h56 : a[0:7] = 8'hAC;
            8'h57 : a[0:7] = 8'hAE;
            8'h58 : a[0:7] = 8'hB0;
            8'h59 : a[0:7] = 8'hB2;
            8'h5A : a[0:7] = 8'hB4;
            8'h5B : a[0:7] = 8'hB6;
            8'h5C : a[0:7] = 8'hB8;
            8'h5D : a[0:7] = 8'hBA;
            8'h5E : a[0:7] = 8'hBC;
            8'h5F : a[0:7] = 8'hBE;
            8'h60 : a[0:7] = 8'hC0;
            8'h61 : a[0:7] = 8'hC2;
            8'h62 : a[0:7] = 8'hC4;
            8'h63 : a[0:7] = 8'hC6;
            8'h64 : a[0:7] = 8'hC8;
            8'h65 : a[0:7] = 8'hCA;
            8'h66 : a[0:7] = 8'hCC;
            8'h67 : a[0:7] = 8'hCE;
            8'h68 : a[0:7] = 8'hD0;
            8'h69 : a[0:7] = 8'hD2;
            8'h6A : a[0:7] = 8'hD4;
            8'h6B : a[0:7] = 8'hD6;
            8'h6C : a[0:7] = 8'hD8;
            8'h6D : a[0:7] = 8'hDA;
            8'h6E : a[0:7] = 8'hDC;
            8'h6F : a[0:7] = 8'hDE;
            8'h70 : a[0:7] = 8'hE0;
            8'h71 : a[0:7] = 8'hE2;
            8'h72 : a[0:7] = 8'hE4;
            8'h73 : a[0:7] = 8'hE6;
            8'h74 : a[0:7] = 8'hE8;
            8'h75 : a[0:7] = 8'hEA;
            8'h76 : a[0:7] = 8'hEC;
            8'h77 : a[0:7] = 8'hEE;
            8'h78 : a[0:7] = 8'hF0;
            8'h79 : a[0:7] = 8'hF2;
            8'h7A : a[0:7] = 8'hF4;
            8'h7B : a[0:7] = 8'hF6;
            8'h7C : a[0:7] = 8'hF8;
            8'h7D : a[0:7] = 8'hFA;
            8'h7E : a[0:7] = 8'hFC;
            8'h7F : a[0:7] = 8'hFE;
            8'h80 : a[0:7] = 8'h1B;
            8'h81 : a[0:7] = 8'h19;
            8'h82 : a[0:7] = 8'h1F;
            8'h83 : a[0:7] = 8'h1D;
            8'h84 : a[0:7] = 8'h13;
            8'h85 : a[0:7] = 8'h11;
            8'h86 : a[0:7] = 8'h17;
            8'h87 : a[0:7] = 8'h15;
            8'h88 : a[0:7] = 8'hB;
            8'h89 : a[0:7] = 8'h9;
            8'h8A : a[0:7] = 8'hF;
            8'h8B : a[0:7] = 8'hD;
            8'h8C : a[0:7] = 8'h3;
            8'h8D : a[0:7] = 8'h1;
            8'h8E : a[0:7] = 8'h7;
            8'h8F : a[0:7] = 8'h5;
            8'h90 : a[0:7] = 8'h3B;
            8'h91 : a[0:7] = 8'h39;
            8'h92 : a[0:7] = 8'h3F;
            8'h93 : a[0:7] = 8'h3D;
            8'h94 : a[0:7] = 8'h33;
            8'h95 : a[0:7] = 8'h31;
            8'h96 : a[0:7] = 8'h37;
            8'h97 : a[0:7] = 8'h35;
            8'h98 : a[0:7] = 8'h2B;
            8'h99 : a[0:7] = 8'h29;
            8'h9A : a[0:7] = 8'h2F;
            8'h9B : a[0:7] = 8'h2D;
            8'h9C : a[0:7] = 8'h23;
            8'h9D : a[0:7] = 8'h21;
            8'h9E : a[0:7] = 8'h27;
            8'h9F : a[0:7] = 8'h25;
            8'hA0 : a[0:7] = 8'h5B;
            8'hA1 : a[0:7] = 8'h59;
            8'hA2 : a[0:7] = 8'h5F;
            8'hA3 : a[0:7] = 8'h5D;
            8'hA4 : a[0:7] = 8'h53;
            8'hA5 : a[0:7] = 8'h51;
            8'hA6 : a[0:7] = 8'h57;
            8'hA7 : a[0:7] = 8'h55;
            8'hA8 : a[0:7] = 8'h4B;
            8'hA9 : a[0:7] = 8'h49;
            8'hAA : a[0:7] = 8'h4F;
            8'hAB : a[0:7] = 8'h4D;
            8'hAC : a[0:7] = 8'h43;
            8'hAD : a[0:7] = 8'h41;
            8'hAE : a[0:7] = 8'h47;
            8'hAF : a[0:7] = 8'h45;
            8'hB0 : a[0:7] = 8'h7B;
            8'hB1 : a[0:7] = 8'h79;
            8'hB2 : a[0:7] = 8'h7F;
            8'hB3 : a[0:7] = 8'h7D;
            8'hB4 : a[0:7] = 8'h73;
            8'hB5 : a[0:7] = 8'h71;
            8'hB6 : a[0:7] = 8'h77;
            8'hB7 : a[0:7] = 8'h75;
            8'hB8 : a[0:7] = 8'h6B;
            8'hB9 : a[0:7] = 8'h69;
            8'hBA : a[0:7] = 8'h6F;
            8'hBB : a[0:7] = 8'h6D;
            8'hBC : a[0:7] = 8'h63;
            8'hBD : a[0:7] = 8'h61;
            8'hBE : a[0:7] = 8'h67;
            8'hBF : a[0:7] = 8'h65;
            8'hC0 : a[0:7] = 8'h9B;
            8'hC1 : a[0:7] = 8'h99;
            8'hC2 : a[0:7] = 8'h9F;
            8'hC3 : a[0:7] = 8'h9D;
            8'hC4 : a[0:7] = 8'h93;
            8'hC5 : a[0:7] = 8'h91;
            8'hC6 : a[0:7] = 8'h97;
            8'hC7 : a[0:7] = 8'h95;
            8'hC8 : a[0:7] = 8'h8B;
            8'hC9 : a[0:7] = 8'h89;
            8'hCA : a[0:7] = 8'h8F;
            8'hCB : a[0:7] = 8'h8D;
            8'hCC : a[0:7] = 8'h83;
            8'hCD : a[0:7] = 8'h81;
            8'hCE : a[0:7] = 8'h87;
            8'hCF : a[0:7] = 8'h85;
            8'hD0 : a[0:7] = 8'hBB;
            8'hD1 : a[0:7] = 8'hB9;
            8'hD2 : a[0:7] = 8'hBF;
            8'hD3 : a[0:7] = 8'hBD;
            8'hD4 : a[0:7] = 8'hB3;
            8'hD5 : a[0:7] = 8'hB1;
            8'hD6 : a[0:7] = 8'hB7;
            8'hD7 : a[0:7] = 8'hB5;
            8'hD8 : a[0:7] = 8'hAB;
            8'hD9 : a[0:7] = 8'hA9;
            8'hDA : a[0:7] = 8'hAF;
            8'hDB : a[0:7] = 8'hAD;
            8'hDC : a[0:7] = 8'hA3;
            8'hDD : a[0:7] = 8'hA1;
            8'hDE : a[0:7] = 8'hA7;
            8'hDF : a[0:7] = 8'hA5;
            8'hE0 : a[0:7] = 8'hDB;
            8'hE1 : a[0:7] = 8'hD9;
            8'hE2 : a[0:7] = 8'hDF;
            8'hE3 : a[0:7] = 8'hDD;
            8'hE4 : a[0:7] = 8'hD3;
            8'hE5 : a[0:7] = 8'hD1;
            8'hE6 : a[0:7] = 8'hD7;
            8'hE7 : a[0:7] = 8'hD5;
            8'hE8 : a[0:7] = 8'hCB;
            8'hE9 : a[0:7] = 8'hC9;
            8'hEA : a[0:7] = 8'hCF;
            8'hEB : a[0:7] = 8'hCD;
            8'hEC : a[0:7] = 8'hC3;
            8'hED : a[0:7] = 8'hC1;
            8'hEE : a[0:7] = 8'hC7;
            8'hEF : a[0:7] = 8'hC5;
            8'hF0 : a[0:7] = 8'hFB;
            8'hF1 : a[0:7] = 8'hF9;
            8'hF2 : a[0:7] = 8'hFF;
            8'hF3 : a[0:7] = 8'hFD;
            8'hF4 : a[0:7] = 8'hF3;
            8'hF5 : a[0:7] = 8'hF1;
            8'hF6 : a[0:7] = 8'hF7;
            8'hF7 : a[0:7] = 8'hF5;
            8'hF8 : a[0:7] = 8'hEB;
            8'hF9 : a[0:7] = 8'hE9;
            8'hFA : a[0:7] = 8'hEF;
            8'hFB : a[0:7] = 8'hED;
            8'hFC : a[0:7] = 8'hE3;
            8'hFD : a[0:7] = 8'hE1;
            8'hFE : a[0:7] = 8'hE7;
            8'hFF : a[0:7] = 8'hE5;
        endcase
    end

    always @(row[8:15]) begin
        // Multiplication with 3
        case (row[8:15])
            8'h0 : b[0:7] = 8'h0;
            8'h1 : b[0:7] = 8'h3;
            8'h2 : b[0:7] = 8'h6;
            8'h3 : b[0:7] = 8'h5;
            8'h4 : b[0:7] = 8'hC;
            8'h5 : b[0:7] = 8'hF;
            8'h6 : b[0:7] = 8'hA;
            8'h7 : b[0:7] = 8'h9;
            8'h8 : b[0:7] = 8'h18;
            8'h9 : b[0:7] = 8'h1B;
            8'hA : b[0:7] = 8'h1E;
            8'hB : b[0:7] = 8'h1D;
            8'hC : b[0:7] = 8'h14;
            8'hD : b[0:7] = 8'h17;
            8'hE : b[0:7] = 8'h12;
            8'hF : b[0:7] = 8'h11;
            8'h10 : b[0:7] = 8'h30;
            8'h11 : b[0:7] = 8'h33;
            8'h12 : b[0:7] = 8'h36;
            8'h13 : b[0:7] = 8'h35;
            8'h14 : b[0:7] = 8'h3C;
            8'h15 : b[0:7] = 8'h3F;
            8'h16 : b[0:7] = 8'h3A;
            8'h17 : b[0:7] = 8'h39;
            8'h18 : b[0:7] = 8'h28;
            8'h19 : b[0:7] = 8'h2B;
            8'h1A : b[0:7] = 8'h2E;
            8'h1B : b[0:7] = 8'h2D;
            8'h1C : b[0:7] = 8'h24;
            8'h1D : b[0:7] = 8'h27;
            8'h1E : b[0:7] = 8'h22;
            8'h1F : b[0:7] = 8'h21;
            8'h20 : b[0:7] = 8'h60;
            8'h21 : b[0:7] = 8'h63;
            8'h22 : b[0:7] = 8'h66;
            8'h23 : b[0:7] = 8'h65;
            8'h24 : b[0:7] = 8'h6C;
            8'h25 : b[0:7] = 8'h6F;
            8'h26 : b[0:7] = 8'h6A;
            8'h27 : b[0:7] = 8'h69;
            8'h28 : b[0:7] = 8'h78;
            8'h29 : b[0:7] = 8'h7B;
            8'h2A : b[0:7] = 8'h7E;
            8'h2B : b[0:7] = 8'h7D;
            8'h2C : b[0:7] = 8'h74;
            8'h2D : b[0:7] = 8'h77;
            8'h2E : b[0:7] = 8'h72;
            8'h2F : b[0:7] = 8'h71;
            8'h30 : b[0:7] = 8'h50;
            8'h31 : b[0:7] = 8'h53;
            8'h32 : b[0:7] = 8'h56;
            8'h33 : b[0:7] = 8'h55;
            8'h34 : b[0:7] = 8'h5C;
            8'h35 : b[0:7] = 8'h5F;
            8'h36 : b[0:7] = 8'h5A;
            8'h37 : b[0:7] = 8'h59;
            8'h38 : b[0:7] = 8'h48;
            8'h39 : b[0:7] = 8'h4B;
            8'h3A : b[0:7] = 8'h4E;
            8'h3B : b[0:7] = 8'h4D;
            8'h3C : b[0:7] = 8'h44;
            8'h3D : b[0:7] = 8'h47;
            8'h3E : b[0:7] = 8'h42;
            8'h3F : b[0:7] = 8'h41;
            8'h40 : b[0:7] = 8'hC0;
            8'h41 : b[0:7] = 8'hC3;
            8'h42 : b[0:7] = 8'hC6;
            8'h43 : b[0:7] = 8'hC5;
            8'h44 : b[0:7] = 8'hCC;
            8'h45 : b[0:7] = 8'hCF;
            8'h46 : b[0:7] = 8'hCA;
            8'h47 : b[0:7] = 8'hC9;
            8'h48 : b[0:7] = 8'hD8;
            8'h49 : b[0:7] = 8'hDB;
            8'h4A : b[0:7] = 8'hDE;
            8'h4B : b[0:7] = 8'hDD;
            8'h4C : b[0:7] = 8'hD4;
            8'h4D : b[0:7] = 8'hD7;
            8'h4E : b[0:7] = 8'hD2;
            8'h4F : b[0:7] = 8'hD1;
            8'h50 : b[0:7] = 8'hF0;
            8'h51 : b[0:7] = 8'hF3;
            8'h52 : b[0:7] = 8'hF6;
            8'h53 : b[0:7] = 8'hF5;
            8'h54 : b[0:7] = 8'hFC;
            8'h55 : b[0:7] = 8'hFF;
            8'h56 : b[0:7] = 8'hFA;
            8'h57 : b[0:7] = 8'hF9;
            8'h58 : b[0:7] = 8'hE8;
            8'h59 : b[0:7] = 8'hEB;
            8'h5A : b[0:7] = 8'hEE;
            8'h5B : b[0:7] = 8'hED;
            8'h5C : b[0:7] = 8'hE4;
            8'h5D : b[0:7] = 8'hE7;
            8'h5E : b[0:7] = 8'hE2;
            8'h5F : b[0:7] = 8'hE1;
            8'h60 : b[0:7] = 8'hA0;
            8'h61 : b[0:7] = 8'hA3;
            8'h62 : b[0:7] = 8'hA6;
            8'h63 : b[0:7] = 8'hA5;
            8'h64 : b[0:7] = 8'hAC;
            8'h65 : b[0:7] = 8'hAF;
            8'h66 : b[0:7] = 8'hAA;
            8'h67 : b[0:7] = 8'hA9;
            8'h68 : b[0:7] = 8'hB8;
            8'h69 : b[0:7] = 8'hBB;
            8'h6A : b[0:7] = 8'hBE;
            8'h6B : b[0:7] = 8'hBD;
            8'h6C : b[0:7] = 8'hB4;
            8'h6D : b[0:7] = 8'hB7;
            8'h6E : b[0:7] = 8'hB2;
            8'h6F : b[0:7] = 8'hB1;
            8'h70 : b[0:7] = 8'h90;
            8'h71 : b[0:7] = 8'h93;
            8'h72 : b[0:7] = 8'h96;
            8'h73 : b[0:7] = 8'h95;
            8'h74 : b[0:7] = 8'h9C;
            8'h75 : b[0:7] = 8'h9F;
            8'h76 : b[0:7] = 8'h9A;
            8'h77 : b[0:7] = 8'h99;
            8'h78 : b[0:7] = 8'h88;
            8'h79 : b[0:7] = 8'h8B;
            8'h7A : b[0:7] = 8'h8E;
            8'h7B : b[0:7] = 8'h8D;
            8'h7C : b[0:7] = 8'h84;
            8'h7D : b[0:7] = 8'h87;
            8'h7E : b[0:7] = 8'h82;
            8'h7F : b[0:7] = 8'h81;
            8'h80 : b[0:7] = 8'h9B;
            8'h81 : b[0:7] = 8'h98;
            8'h82 : b[0:7] = 8'h9D;
            8'h83 : b[0:7] = 8'h9E;
            8'h84 : b[0:7] = 8'h97;
            8'h85 : b[0:7] = 8'h94;
            8'h86 : b[0:7] = 8'h91;
            8'h87 : b[0:7] = 8'h92;
            8'h88 : b[0:7] = 8'h83;
            8'h89 : b[0:7] = 8'h80;
            8'h8A : b[0:7] = 8'h85;
            8'h8B : b[0:7] = 8'h86;
            8'h8C : b[0:7] = 8'h8F;
            8'h8D : b[0:7] = 8'h8C;
            8'h8E : b[0:7] = 8'h89;
            8'h8F : b[0:7] = 8'h8A;
            8'h90 : b[0:7] = 8'hAB;
            8'h91 : b[0:7] = 8'hA8;
            8'h92 : b[0:7] = 8'hAD;
            8'h93 : b[0:7] = 8'hAE;
            8'h94 : b[0:7] = 8'hA7;
            8'h95 : b[0:7] = 8'hA4;
            8'h96 : b[0:7] = 8'hA1;
            8'h97 : b[0:7] = 8'hA2;
            8'h98 : b[0:7] = 8'hB3;
            8'h99 : b[0:7] = 8'hB0;
            8'h9A : b[0:7] = 8'hB5;
            8'h9B : b[0:7] = 8'hB6;
            8'h9C : b[0:7] = 8'hBF;
            8'h9D : b[0:7] = 8'hBC;
            8'h9E : b[0:7] = 8'hB9;
            8'h9F : b[0:7] = 8'hBA;
            8'hA0 : b[0:7] = 8'hFB;
            8'hA1 : b[0:7] = 8'hF8;
            8'hA2 : b[0:7] = 8'hFD;
            8'hA3 : b[0:7] = 8'hFE;
            8'hA4 : b[0:7] = 8'hF7;
            8'hA5 : b[0:7] = 8'hF4;
            8'hA6 : b[0:7] = 8'hF1;
            8'hA7 : b[0:7] = 8'hF2;
            8'hA8 : b[0:7] = 8'hE3;
            8'hA9 : b[0:7] = 8'hE0;
            8'hAA : b[0:7] = 8'hE5;
            8'hAB : b[0:7] = 8'hE6;
            8'hAC : b[0:7] = 8'hEF;
            8'hAD : b[0:7] = 8'hEC;
            8'hAE : b[0:7] = 8'hE9;
            8'hAF : b[0:7] = 8'hEA;
            8'hB0 : b[0:7] = 8'hCB;
            8'hB1 : b[0:7] = 8'hC8;
            8'hB2 : b[0:7] = 8'hCD;
            8'hB3 : b[0:7] = 8'hCE;
            8'hB4 : b[0:7] = 8'hC7;
            8'hB5 : b[0:7] = 8'hC4;
            8'hB6 : b[0:7] = 8'hC1;
            8'hB7 : b[0:7] = 8'hC2;
            8'hB8 : b[0:7] = 8'hD3;
            8'hB9 : b[0:7] = 8'hD0;
            8'hBA : b[0:7] = 8'hD5;
            8'hBB : b[0:7] = 8'hD6;
            8'hBC : b[0:7] = 8'hDF;
            8'hBD : b[0:7] = 8'hDC;
            8'hBE : b[0:7] = 8'hD9;
            8'hBF : b[0:7] = 8'hDA;
            8'hC0 : b[0:7] = 8'h5B;
            8'hC1 : b[0:7] = 8'h58;
            8'hC2 : b[0:7] = 8'h5D;
            8'hC3 : b[0:7] = 8'h5E;
            8'hC4 : b[0:7] = 8'h57;
            8'hC5 : b[0:7] = 8'h54;
            8'hC6 : b[0:7] = 8'h51;
            8'hC7 : b[0:7] = 8'h52;
            8'hC8 : b[0:7] = 8'h43;
            8'hC9 : b[0:7] = 8'h40;
            8'hCA : b[0:7] = 8'h45;
            8'hCB : b[0:7] = 8'h46;
            8'hCC : b[0:7] = 8'h4F;
            8'hCD : b[0:7] = 8'h4C;
            8'hCE : b[0:7] = 8'h49;
            8'hCF : b[0:7] = 8'h4A;
            8'hD0 : b[0:7] = 8'h6B;
            8'hD1 : b[0:7] = 8'h68;
            8'hD2 : b[0:7] = 8'h6D;
            8'hD3 : b[0:7] = 8'h6E;
            8'hD4 : b[0:7] = 8'h67;
            8'hD5 : b[0:7] = 8'h64;
            8'hD6 : b[0:7] = 8'h61;
            8'hD7 : b[0:7] = 8'h62;
            8'hD8 : b[0:7] = 8'h73;
            8'hD9 : b[0:7] = 8'h70;
            8'hDA : b[0:7] = 8'h75;
            8'hDB : b[0:7] = 8'h76;
            8'hDC : b[0:7] = 8'h7F;
            8'hDD : b[0:7] = 8'h7C;
            8'hDE : b[0:7] = 8'h79;
            8'hDF : b[0:7] = 8'h7A;
            8'hE0 : b[0:7] = 8'h3B;
            8'hE1 : b[0:7] = 8'h38;
            8'hE2 : b[0:7] = 8'h3D;
            8'hE3 : b[0:7] = 8'h3E;
            8'hE4 : b[0:7] = 8'h37;
            8'hE5 : b[0:7] = 8'h34;
            8'hE6 : b[0:7] = 8'h31;
            8'hE7 : b[0:7] = 8'h32;
            8'hE8 : b[0:7] = 8'h23;
            8'hE9 : b[0:7] = 8'h20;
            8'hEA : b[0:7] = 8'h25;
            8'hEB : b[0:7] = 8'h26;
            8'hEC : b[0:7] = 8'h2F;
            8'hED : b[0:7] = 8'h2C;
            8'hEE : b[0:7] = 8'h29;
            8'hEF : b[0:7] = 8'h2A;
            8'hF0 : b[0:7] = 8'hB;
            8'hF1 : b[0:7] = 8'h8;
            8'hF2 : b[0:7] = 8'hD;
            8'hF3 : b[0:7] = 8'hE;
            8'hF4 : b[0:7] = 8'h7;
            8'hF5 : b[0:7] = 8'h4;
            8'hF6 : b[0:7] = 8'h1;
            8'hF7 : b[0:7] = 8'h2;
            8'hF8 : b[0:7] = 8'h13;
            8'hF9 : b[0:7] = 8'h10;
            8'hFA : b[0:7] = 8'h15;
            8'hFB : b[0:7] = 8'h16;
            8'hFC : b[0:7] = 8'h1F;
            8'hFD : b[0:7] = 8'h1C;
            8'hFE : b[0:7] = 8'h19;
            8'hFF : b[0:7] = 8'h1A;
        endcase
    end

    // Multiplication with 1
    always @(row[16:23]) begin
        c[0:7] = row[16:23];
    end

    // Multiplication with 1
    always @(row[24:31]) begin
        d[0:7] = row[24:31];
    end

    assign output_row = a ^ b ^ c ^ d;
    
endmodule


module MixColumn2Row (
    input wire [0:31] row,
    output wire [0:7] output_row
);
    reg [0:7] a, b, c, d;

    // Multiplication with 2
    always @(row[8:15]) begin
        case (row[8:15])
            8'h0 : a[0:7] = 8'h0;
            8'h1 : a[0:7] = 8'h2;
            8'h2 : a[0:7] = 8'h4;
            8'h3 : a[0:7] = 8'h6;
            8'h4 : a[0:7] = 8'h8;
            8'h5 : a[0:7] = 8'hA;
            8'h6 : a[0:7] = 8'hC;
            8'h7 : a[0:7] = 8'hE;
            8'h8 : a[0:7] = 8'h10;
            8'h9 : a[0:7] = 8'h12;
            8'hA : a[0:7] = 8'h14;
            8'hB : a[0:7] = 8'h16;
            8'hC : a[0:7] = 8'h18;
            8'hD : a[0:7] = 8'h1A;
            8'hE : a[0:7] = 8'h1C;
            8'hF : a[0:7] = 8'h1E;
            8'h10 : a[0:7] = 8'h20;
            8'h11 : a[0:7] = 8'h22;
            8'h12 : a[0:7] = 8'h24;
            8'h13 : a[0:7] = 8'h26;
            8'h14 : a[0:7] = 8'h28;
            8'h15 : a[0:7] = 8'h2A;
            8'h16 : a[0:7] = 8'h2C;
            8'h17 : a[0:7] = 8'h2E;
            8'h18 : a[0:7] = 8'h30;
            8'h19 : a[0:7] = 8'h32;
            8'h1A : a[0:7] = 8'h34;
            8'h1B : a[0:7] = 8'h36;
            8'h1C : a[0:7] = 8'h38;
            8'h1D : a[0:7] = 8'h3A;
            8'h1E : a[0:7] = 8'h3C;
            8'h1F : a[0:7] = 8'h3E;
            8'h20 : a[0:7] = 8'h40;
            8'h21 : a[0:7] = 8'h42;
            8'h22 : a[0:7] = 8'h44;
            8'h23 : a[0:7] = 8'h46;
            8'h24 : a[0:7] = 8'h48;
            8'h25 : a[0:7] = 8'h4A;
            8'h26 : a[0:7] = 8'h4C;
            8'h27 : a[0:7] = 8'h4E;
            8'h28 : a[0:7] = 8'h50;
            8'h29 : a[0:7] = 8'h52;
            8'h2A : a[0:7] = 8'h54;
            8'h2B : a[0:7] = 8'h56;
            8'h2C : a[0:7] = 8'h58;
            8'h2D : a[0:7] = 8'h5A;
            8'h2E : a[0:7] = 8'h5C;
            8'h2F : a[0:7] = 8'h5E;
            8'h30 : a[0:7] = 8'h60;
            8'h31 : a[0:7] = 8'h62;
            8'h32 : a[0:7] = 8'h64;
            8'h33 : a[0:7] = 8'h66;
            8'h34 : a[0:7] = 8'h68;
            8'h35 : a[0:7] = 8'h6A;
            8'h36 : a[0:7] = 8'h6C;
            8'h37 : a[0:7] = 8'h6E;
            8'h38 : a[0:7] = 8'h70;
            8'h39 : a[0:7] = 8'h72;
            8'h3A : a[0:7] = 8'h74;
            8'h3B : a[0:7] = 8'h76;
            8'h3C : a[0:7] = 8'h78;
            8'h3D : a[0:7] = 8'h7A;
            8'h3E : a[0:7] = 8'h7C;
            8'h3F : a[0:7] = 8'h7E;
            8'h40 : a[0:7] = 8'h80;
            8'h41 : a[0:7] = 8'h82;
            8'h42 : a[0:7] = 8'h84;
            8'h43 : a[0:7] = 8'h86;
            8'h44 : a[0:7] = 8'h88;
            8'h45 : a[0:7] = 8'h8A;
            8'h46 : a[0:7] = 8'h8C;
            8'h47 : a[0:7] = 8'h8E;
            8'h48 : a[0:7] = 8'h90;
            8'h49 : a[0:7] = 8'h92;
            8'h4A : a[0:7] = 8'h94;
            8'h4B : a[0:7] = 8'h96;
            8'h4C : a[0:7] = 8'h98;
            8'h4D : a[0:7] = 8'h9A;
            8'h4E : a[0:7] = 8'h9C;
            8'h4F : a[0:7] = 8'h9E;
            8'h50 : a[0:7] = 8'hA0;
            8'h51 : a[0:7] = 8'hA2;
            8'h52 : a[0:7] = 8'hA4;
            8'h53 : a[0:7] = 8'hA6;
            8'h54 : a[0:7] = 8'hA8;
            8'h55 : a[0:7] = 8'hAA;
            8'h56 : a[0:7] = 8'hAC;
            8'h57 : a[0:7] = 8'hAE;
            8'h58 : a[0:7] = 8'hB0;
            8'h59 : a[0:7] = 8'hB2;
            8'h5A : a[0:7] = 8'hB4;
            8'h5B : a[0:7] = 8'hB6;
            8'h5C : a[0:7] = 8'hB8;
            8'h5D : a[0:7] = 8'hBA;
            8'h5E : a[0:7] = 8'hBC;
            8'h5F : a[0:7] = 8'hBE;
            8'h60 : a[0:7] = 8'hC0;
            8'h61 : a[0:7] = 8'hC2;
            8'h62 : a[0:7] = 8'hC4;
            8'h63 : a[0:7] = 8'hC6;
            8'h64 : a[0:7] = 8'hC8;
            8'h65 : a[0:7] = 8'hCA;
            8'h66 : a[0:7] = 8'hCC;
            8'h67 : a[0:7] = 8'hCE;
            8'h68 : a[0:7] = 8'hD0;
            8'h69 : a[0:7] = 8'hD2;
            8'h6A : a[0:7] = 8'hD4;
            8'h6B : a[0:7] = 8'hD6;
            8'h6C : a[0:7] = 8'hD8;
            8'h6D : a[0:7] = 8'hDA;
            8'h6E : a[0:7] = 8'hDC;
            8'h6F : a[0:7] = 8'hDE;
            8'h70 : a[0:7] = 8'hE0;
            8'h71 : a[0:7] = 8'hE2;
            8'h72 : a[0:7] = 8'hE4;
            8'h73 : a[0:7] = 8'hE6;
            8'h74 : a[0:7] = 8'hE8;
            8'h75 : a[0:7] = 8'hEA;
            8'h76 : a[0:7] = 8'hEC;
            8'h77 : a[0:7] = 8'hEE;
            8'h78 : a[0:7] = 8'hF0;
            8'h79 : a[0:7] = 8'hF2;
            8'h7A : a[0:7] = 8'hF4;
            8'h7B : a[0:7] = 8'hF6;
            8'h7C : a[0:7] = 8'hF8;
            8'h7D : a[0:7] = 8'hFA;
            8'h7E : a[0:7] = 8'hFC;
            8'h7F : a[0:7] = 8'hFE;
            8'h80 : a[0:7] = 8'h1B;
            8'h81 : a[0:7] = 8'h19;
            8'h82 : a[0:7] = 8'h1F;
            8'h83 : a[0:7] = 8'h1D;
            8'h84 : a[0:7] = 8'h13;
            8'h85 : a[0:7] = 8'h11;
            8'h86 : a[0:7] = 8'h17;
            8'h87 : a[0:7] = 8'h15;
            8'h88 : a[0:7] = 8'hB;
            8'h89 : a[0:7] = 8'h9;
            8'h8A : a[0:7] = 8'hF;
            8'h8B : a[0:7] = 8'hD;
            8'h8C : a[0:7] = 8'h3;
            8'h8D : a[0:7] = 8'h1;
            8'h8E : a[0:7] = 8'h7;
            8'h8F : a[0:7] = 8'h5;
            8'h90 : a[0:7] = 8'h3B;
            8'h91 : a[0:7] = 8'h39;
            8'h92 : a[0:7] = 8'h3F;
            8'h93 : a[0:7] = 8'h3D;
            8'h94 : a[0:7] = 8'h33;
            8'h95 : a[0:7] = 8'h31;
            8'h96 : a[0:7] = 8'h37;
            8'h97 : a[0:7] = 8'h35;
            8'h98 : a[0:7] = 8'h2B;
            8'h99 : a[0:7] = 8'h29;
            8'h9A : a[0:7] = 8'h2F;
            8'h9B : a[0:7] = 8'h2D;
            8'h9C : a[0:7] = 8'h23;
            8'h9D : a[0:7] = 8'h21;
            8'h9E : a[0:7] = 8'h27;
            8'h9F : a[0:7] = 8'h25;
            8'hA0 : a[0:7] = 8'h5B;
            8'hA1 : a[0:7] = 8'h59;
            8'hA2 : a[0:7] = 8'h5F;
            8'hA3 : a[0:7] = 8'h5D;
            8'hA4 : a[0:7] = 8'h53;
            8'hA5 : a[0:7] = 8'h51;
            8'hA6 : a[0:7] = 8'h57;
            8'hA7 : a[0:7] = 8'h55;
            8'hA8 : a[0:7] = 8'h4B;
            8'hA9 : a[0:7] = 8'h49;
            8'hAA : a[0:7] = 8'h4F;
            8'hAB : a[0:7] = 8'h4D;
            8'hAC : a[0:7] = 8'h43;
            8'hAD : a[0:7] = 8'h41;
            8'hAE : a[0:7] = 8'h47;
            8'hAF : a[0:7] = 8'h45;
            8'hB0 : a[0:7] = 8'h7B;
            8'hB1 : a[0:7] = 8'h79;
            8'hB2 : a[0:7] = 8'h7F;
            8'hB3 : a[0:7] = 8'h7D;
            8'hB4 : a[0:7] = 8'h73;
            8'hB5 : a[0:7] = 8'h71;
            8'hB6 : a[0:7] = 8'h77;
            8'hB7 : a[0:7] = 8'h75;
            8'hB8 : a[0:7] = 8'h6B;
            8'hB9 : a[0:7] = 8'h69;
            8'hBA : a[0:7] = 8'h6F;
            8'hBB : a[0:7] = 8'h6D;
            8'hBC : a[0:7] = 8'h63;
            8'hBD : a[0:7] = 8'h61;
            8'hBE : a[0:7] = 8'h67;
            8'hBF : a[0:7] = 8'h65;
            8'hC0 : a[0:7] = 8'h9B;
            8'hC1 : a[0:7] = 8'h99;
            8'hC2 : a[0:7] = 8'h9F;
            8'hC3 : a[0:7] = 8'h9D;
            8'hC4 : a[0:7] = 8'h93;
            8'hC5 : a[0:7] = 8'h91;
            8'hC6 : a[0:7] = 8'h97;
            8'hC7 : a[0:7] = 8'h95;
            8'hC8 : a[0:7] = 8'h8B;
            8'hC9 : a[0:7] = 8'h89;
            8'hCA : a[0:7] = 8'h8F;
            8'hCB : a[0:7] = 8'h8D;
            8'hCC : a[0:7] = 8'h83;
            8'hCD : a[0:7] = 8'h81;
            8'hCE : a[0:7] = 8'h87;
            8'hCF : a[0:7] = 8'h85;
            8'hD0 : a[0:7] = 8'hBB;
            8'hD1 : a[0:7] = 8'hB9;
            8'hD2 : a[0:7] = 8'hBF;
            8'hD3 : a[0:7] = 8'hBD;
            8'hD4 : a[0:7] = 8'hB3;
            8'hD5 : a[0:7] = 8'hB1;
            8'hD6 : a[0:7] = 8'hB7;
            8'hD7 : a[0:7] = 8'hB5;
            8'hD8 : a[0:7] = 8'hAB;
            8'hD9 : a[0:7] = 8'hA9;
            8'hDA : a[0:7] = 8'hAF;
            8'hDB : a[0:7] = 8'hAD;
            8'hDC : a[0:7] = 8'hA3;
            8'hDD : a[0:7] = 8'hA1;
            8'hDE : a[0:7] = 8'hA7;
            8'hDF : a[0:7] = 8'hA5;
            8'hE0 : a[0:7] = 8'hDB;
            8'hE1 : a[0:7] = 8'hD9;
            8'hE2 : a[0:7] = 8'hDF;
            8'hE3 : a[0:7] = 8'hDD;
            8'hE4 : a[0:7] = 8'hD3;
            8'hE5 : a[0:7] = 8'hD1;
            8'hE6 : a[0:7] = 8'hD7;
            8'hE7 : a[0:7] = 8'hD5;
            8'hE8 : a[0:7] = 8'hCB;
            8'hE9 : a[0:7] = 8'hC9;
            8'hEA : a[0:7] = 8'hCF;
            8'hEB : a[0:7] = 8'hCD;
            8'hEC : a[0:7] = 8'hC3;
            8'hED : a[0:7] = 8'hC1;
            8'hEE : a[0:7] = 8'hC7;
            8'hEF : a[0:7] = 8'hC5;
            8'hF0 : a[0:7] = 8'hFB;
            8'hF1 : a[0:7] = 8'hF9;
            8'hF2 : a[0:7] = 8'hFF;
            8'hF3 : a[0:7] = 8'hFD;
            8'hF4 : a[0:7] = 8'hF3;
            8'hF5 : a[0:7] = 8'hF1;
            8'hF6 : a[0:7] = 8'hF7;
            8'hF7 : a[0:7] = 8'hF5;
            8'hF8 : a[0:7] = 8'hEB;
            8'hF9 : a[0:7] = 8'hE9;
            8'hFA : a[0:7] = 8'hEF;
            8'hFB : a[0:7] = 8'hED;
            8'hFC : a[0:7] = 8'hE3;
            8'hFD : a[0:7] = 8'hE1;
            8'hFE : a[0:7] = 8'hE7;
            8'hFF : a[0:7] = 8'hE5;
        endcase
    end

    always @(row[16:23]) begin
        // Multiplication with 3
        case (row[16:23])
            8'h0 : b[0:7] = 8'h0;
            8'h1 : b[0:7] = 8'h3;
            8'h2 : b[0:7] = 8'h6;
            8'h3 : b[0:7] = 8'h5;
            8'h4 : b[0:7] = 8'hC;
            8'h5 : b[0:7] = 8'hF;
            8'h6 : b[0:7] = 8'hA;
            8'h7 : b[0:7] = 8'h9;
            8'h8 : b[0:7] = 8'h18;
            8'h9 : b[0:7] = 8'h1B;
            8'hA : b[0:7] = 8'h1E;
            8'hB : b[0:7] = 8'h1D;
            8'hC : b[0:7] = 8'h14;
            8'hD : b[0:7] = 8'h17;
            8'hE : b[0:7] = 8'h12;
            8'hF : b[0:7] = 8'h11;
            8'h10 : b[0:7] = 8'h30;
            8'h11 : b[0:7] = 8'h33;
            8'h12 : b[0:7] = 8'h36;
            8'h13 : b[0:7] = 8'h35;
            8'h14 : b[0:7] = 8'h3C;
            8'h15 : b[0:7] = 8'h3F;
            8'h16 : b[0:7] = 8'h3A;
            8'h17 : b[0:7] = 8'h39;
            8'h18 : b[0:7] = 8'h28;
            8'h19 : b[0:7] = 8'h2B;
            8'h1A : b[0:7] = 8'h2E;
            8'h1B : b[0:7] = 8'h2D;
            8'h1C : b[0:7] = 8'h24;
            8'h1D : b[0:7] = 8'h27;
            8'h1E : b[0:7] = 8'h22;
            8'h1F : b[0:7] = 8'h21;
            8'h20 : b[0:7] = 8'h60;
            8'h21 : b[0:7] = 8'h63;
            8'h22 : b[0:7] = 8'h66;
            8'h23 : b[0:7] = 8'h65;
            8'h24 : b[0:7] = 8'h6C;
            8'h25 : b[0:7] = 8'h6F;
            8'h26 : b[0:7] = 8'h6A;
            8'h27 : b[0:7] = 8'h69;
            8'h28 : b[0:7] = 8'h78;
            8'h29 : b[0:7] = 8'h7B;
            8'h2A : b[0:7] = 8'h7E;
            8'h2B : b[0:7] = 8'h7D;
            8'h2C : b[0:7] = 8'h74;
            8'h2D : b[0:7] = 8'h77;
            8'h2E : b[0:7] = 8'h72;
            8'h2F : b[0:7] = 8'h71;
            8'h30 : b[0:7] = 8'h50;
            8'h31 : b[0:7] = 8'h53;
            8'h32 : b[0:7] = 8'h56;
            8'h33 : b[0:7] = 8'h55;
            8'h34 : b[0:7] = 8'h5C;
            8'h35 : b[0:7] = 8'h5F;
            8'h36 : b[0:7] = 8'h5A;
            8'h37 : b[0:7] = 8'h59;
            8'h38 : b[0:7] = 8'h48;
            8'h39 : b[0:7] = 8'h4B;
            8'h3A : b[0:7] = 8'h4E;
            8'h3B : b[0:7] = 8'h4D;
            8'h3C : b[0:7] = 8'h44;
            8'h3D : b[0:7] = 8'h47;
            8'h3E : b[0:7] = 8'h42;
            8'h3F : b[0:7] = 8'h41;
            8'h40 : b[0:7] = 8'hC0;
            8'h41 : b[0:7] = 8'hC3;
            8'h42 : b[0:7] = 8'hC6;
            8'h43 : b[0:7] = 8'hC5;
            8'h44 : b[0:7] = 8'hCC;
            8'h45 : b[0:7] = 8'hCF;
            8'h46 : b[0:7] = 8'hCA;
            8'h47 : b[0:7] = 8'hC9;
            8'h48 : b[0:7] = 8'hD8;
            8'h49 : b[0:7] = 8'hDB;
            8'h4A : b[0:7] = 8'hDE;
            8'h4B : b[0:7] = 8'hDD;
            8'h4C : b[0:7] = 8'hD4;
            8'h4D : b[0:7] = 8'hD7;
            8'h4E : b[0:7] = 8'hD2;
            8'h4F : b[0:7] = 8'hD1;
            8'h50 : b[0:7] = 8'hF0;
            8'h51 : b[0:7] = 8'hF3;
            8'h52 : b[0:7] = 8'hF6;
            8'h53 : b[0:7] = 8'hF5;
            8'h54 : b[0:7] = 8'hFC;
            8'h55 : b[0:7] = 8'hFF;
            8'h56 : b[0:7] = 8'hFA;
            8'h57 : b[0:7] = 8'hF9;
            8'h58 : b[0:7] = 8'hE8;
            8'h59 : b[0:7] = 8'hEB;
            8'h5A : b[0:7] = 8'hEE;
            8'h5B : b[0:7] = 8'hED;
            8'h5C : b[0:7] = 8'hE4;
            8'h5D : b[0:7] = 8'hE7;
            8'h5E : b[0:7] = 8'hE2;
            8'h5F : b[0:7] = 8'hE1;
            8'h60 : b[0:7] = 8'hA0;
            8'h61 : b[0:7] = 8'hA3;
            8'h62 : b[0:7] = 8'hA6;
            8'h63 : b[0:7] = 8'hA5;
            8'h64 : b[0:7] = 8'hAC;
            8'h65 : b[0:7] = 8'hAF;
            8'h66 : b[0:7] = 8'hAA;
            8'h67 : b[0:7] = 8'hA9;
            8'h68 : b[0:7] = 8'hB8;
            8'h69 : b[0:7] = 8'hBB;
            8'h6A : b[0:7] = 8'hBE;
            8'h6B : b[0:7] = 8'hBD;
            8'h6C : b[0:7] = 8'hB4;
            8'h6D : b[0:7] = 8'hB7;
            8'h6E : b[0:7] = 8'hB2;
            8'h6F : b[0:7] = 8'hB1;
            8'h70 : b[0:7] = 8'h90;
            8'h71 : b[0:7] = 8'h93;
            8'h72 : b[0:7] = 8'h96;
            8'h73 : b[0:7] = 8'h95;
            8'h74 : b[0:7] = 8'h9C;
            8'h75 : b[0:7] = 8'h9F;
            8'h76 : b[0:7] = 8'h9A;
            8'h77 : b[0:7] = 8'h99;
            8'h78 : b[0:7] = 8'h88;
            8'h79 : b[0:7] = 8'h8B;
            8'h7A : b[0:7] = 8'h8E;
            8'h7B : b[0:7] = 8'h8D;
            8'h7C : b[0:7] = 8'h84;
            8'h7D : b[0:7] = 8'h87;
            8'h7E : b[0:7] = 8'h82;
            8'h7F : b[0:7] = 8'h81;
            8'h80 : b[0:7] = 8'h9B;
            8'h81 : b[0:7] = 8'h98;
            8'h82 : b[0:7] = 8'h9D;
            8'h83 : b[0:7] = 8'h9E;
            8'h84 : b[0:7] = 8'h97;
            8'h85 : b[0:7] = 8'h94;
            8'h86 : b[0:7] = 8'h91;
            8'h87 : b[0:7] = 8'h92;
            8'h88 : b[0:7] = 8'h83;
            8'h89 : b[0:7] = 8'h80;
            8'h8A : b[0:7] = 8'h85;
            8'h8B : b[0:7] = 8'h86;
            8'h8C : b[0:7] = 8'h8F;
            8'h8D : b[0:7] = 8'h8C;
            8'h8E : b[0:7] = 8'h89;
            8'h8F : b[0:7] = 8'h8A;
            8'h90 : b[0:7] = 8'hAB;
            8'h91 : b[0:7] = 8'hA8;
            8'h92 : b[0:7] = 8'hAD;
            8'h93 : b[0:7] = 8'hAE;
            8'h94 : b[0:7] = 8'hA7;
            8'h95 : b[0:7] = 8'hA4;
            8'h96 : b[0:7] = 8'hA1;
            8'h97 : b[0:7] = 8'hA2;
            8'h98 : b[0:7] = 8'hB3;
            8'h99 : b[0:7] = 8'hB0;
            8'h9A : b[0:7] = 8'hB5;
            8'h9B : b[0:7] = 8'hB6;
            8'h9C : b[0:7] = 8'hBF;
            8'h9D : b[0:7] = 8'hBC;
            8'h9E : b[0:7] = 8'hB9;
            8'h9F : b[0:7] = 8'hBA;
            8'hA0 : b[0:7] = 8'hFB;
            8'hA1 : b[0:7] = 8'hF8;
            8'hA2 : b[0:7] = 8'hFD;
            8'hA3 : b[0:7] = 8'hFE;
            8'hA4 : b[0:7] = 8'hF7;
            8'hA5 : b[0:7] = 8'hF4;
            8'hA6 : b[0:7] = 8'hF1;
            8'hA7 : b[0:7] = 8'hF2;
            8'hA8 : b[0:7] = 8'hE3;
            8'hA9 : b[0:7] = 8'hE0;
            8'hAA : b[0:7] = 8'hE5;
            8'hAB : b[0:7] = 8'hE6;
            8'hAC : b[0:7] = 8'hEF;
            8'hAD : b[0:7] = 8'hEC;
            8'hAE : b[0:7] = 8'hE9;
            8'hAF : b[0:7] = 8'hEA;
            8'hB0 : b[0:7] = 8'hCB;
            8'hB1 : b[0:7] = 8'hC8;
            8'hB2 : b[0:7] = 8'hCD;
            8'hB3 : b[0:7] = 8'hCE;
            8'hB4 : b[0:7] = 8'hC7;
            8'hB5 : b[0:7] = 8'hC4;
            8'hB6 : b[0:7] = 8'hC1;
            8'hB7 : b[0:7] = 8'hC2;
            8'hB8 : b[0:7] = 8'hD3;
            8'hB9 : b[0:7] = 8'hD0;
            8'hBA : b[0:7] = 8'hD5;
            8'hBB : b[0:7] = 8'hD6;
            8'hBC : b[0:7] = 8'hDF;
            8'hBD : b[0:7] = 8'hDC;
            8'hBE : b[0:7] = 8'hD9;
            8'hBF : b[0:7] = 8'hDA;
            8'hC0 : b[0:7] = 8'h5B;
            8'hC1 : b[0:7] = 8'h58;
            8'hC2 : b[0:7] = 8'h5D;
            8'hC3 : b[0:7] = 8'h5E;
            8'hC4 : b[0:7] = 8'h57;
            8'hC5 : b[0:7] = 8'h54;
            8'hC6 : b[0:7] = 8'h51;
            8'hC7 : b[0:7] = 8'h52;
            8'hC8 : b[0:7] = 8'h43;
            8'hC9 : b[0:7] = 8'h40;
            8'hCA : b[0:7] = 8'h45;
            8'hCB : b[0:7] = 8'h46;
            8'hCC : b[0:7] = 8'h4F;
            8'hCD : b[0:7] = 8'h4C;
            8'hCE : b[0:7] = 8'h49;
            8'hCF : b[0:7] = 8'h4A;
            8'hD0 : b[0:7] = 8'h6B;
            8'hD1 : b[0:7] = 8'h68;
            8'hD2 : b[0:7] = 8'h6D;
            8'hD3 : b[0:7] = 8'h6E;
            8'hD4 : b[0:7] = 8'h67;
            8'hD5 : b[0:7] = 8'h64;
            8'hD6 : b[0:7] = 8'h61;
            8'hD7 : b[0:7] = 8'h62;
            8'hD8 : b[0:7] = 8'h73;
            8'hD9 : b[0:7] = 8'h70;
            8'hDA : b[0:7] = 8'h75;
            8'hDB : b[0:7] = 8'h76;
            8'hDC : b[0:7] = 8'h7F;
            8'hDD : b[0:7] = 8'h7C;
            8'hDE : b[0:7] = 8'h79;
            8'hDF : b[0:7] = 8'h7A;
            8'hE0 : b[0:7] = 8'h3B;
            8'hE1 : b[0:7] = 8'h38;
            8'hE2 : b[0:7] = 8'h3D;
            8'hE3 : b[0:7] = 8'h3E;
            8'hE4 : b[0:7] = 8'h37;
            8'hE5 : b[0:7] = 8'h34;
            8'hE6 : b[0:7] = 8'h31;
            8'hE7 : b[0:7] = 8'h32;
            8'hE8 : b[0:7] = 8'h23;
            8'hE9 : b[0:7] = 8'h20;
            8'hEA : b[0:7] = 8'h25;
            8'hEB : b[0:7] = 8'h26;
            8'hEC : b[0:7] = 8'h2F;
            8'hED : b[0:7] = 8'h2C;
            8'hEE : b[0:7] = 8'h29;
            8'hEF : b[0:7] = 8'h2A;
            8'hF0 : b[0:7] = 8'hB;
            8'hF1 : b[0:7] = 8'h8;
            8'hF2 : b[0:7] = 8'hD;
            8'hF3 : b[0:7] = 8'hE;
            8'hF4 : b[0:7] = 8'h7;
            8'hF5 : b[0:7] = 8'h4;
            8'hF6 : b[0:7] = 8'h1;
            8'hF7 : b[0:7] = 8'h2;
            8'hF8 : b[0:7] = 8'h13;
            8'hF9 : b[0:7] = 8'h10;
            8'hFA : b[0:7] = 8'h15;
            8'hFB : b[0:7] = 8'h16;
            8'hFC : b[0:7] = 8'h1F;
            8'hFD : b[0:7] = 8'h1C;
            8'hFE : b[0:7] = 8'h19;
            8'hFF : b[0:7] = 8'h1A;
        endcase
    end

    // Multiplication with 1
    always @(row[0:7]) begin
        c[0:7] = row[0:7];
    end

    // Multiplication with 1
    always @(row[24:31]) begin
        d[0:7] = row[24:31];
    end

    assign output_row = a ^ b ^ c ^ d;
    
endmodule


module MixColumn3Row (
    input wire [0:31] row,
    output wire [0:7] output_row
);
    reg [0:7] a, b, c, d;

    // Multiplication with 2
    always @(row[16:23]) begin
        case (row[16:23])
            8'h0 : a[0:7] = 8'h0;
            8'h1 : a[0:7] = 8'h2;
            8'h2 : a[0:7] = 8'h4;
            8'h3 : a[0:7] = 8'h6;
            8'h4 : a[0:7] = 8'h8;
            8'h5 : a[0:7] = 8'hA;
            8'h6 : a[0:7] = 8'hC;
            8'h7 : a[0:7] = 8'hE;
            8'h8 : a[0:7] = 8'h10;
            8'h9 : a[0:7] = 8'h12;
            8'hA : a[0:7] = 8'h14;
            8'hB : a[0:7] = 8'h16;
            8'hC : a[0:7] = 8'h18;
            8'hD : a[0:7] = 8'h1A;
            8'hE : a[0:7] = 8'h1C;
            8'hF : a[0:7] = 8'h1E;
            8'h10 : a[0:7] = 8'h20;
            8'h11 : a[0:7] = 8'h22;
            8'h12 : a[0:7] = 8'h24;
            8'h13 : a[0:7] = 8'h26;
            8'h14 : a[0:7] = 8'h28;
            8'h15 : a[0:7] = 8'h2A;
            8'h16 : a[0:7] = 8'h2C;
            8'h17 : a[0:7] = 8'h2E;
            8'h18 : a[0:7] = 8'h30;
            8'h19 : a[0:7] = 8'h32;
            8'h1A : a[0:7] = 8'h34;
            8'h1B : a[0:7] = 8'h36;
            8'h1C : a[0:7] = 8'h38;
            8'h1D : a[0:7] = 8'h3A;
            8'h1E : a[0:7] = 8'h3C;
            8'h1F : a[0:7] = 8'h3E;
            8'h20 : a[0:7] = 8'h40;
            8'h21 : a[0:7] = 8'h42;
            8'h22 : a[0:7] = 8'h44;
            8'h23 : a[0:7] = 8'h46;
            8'h24 : a[0:7] = 8'h48;
            8'h25 : a[0:7] = 8'h4A;
            8'h26 : a[0:7] = 8'h4C;
            8'h27 : a[0:7] = 8'h4E;
            8'h28 : a[0:7] = 8'h50;
            8'h29 : a[0:7] = 8'h52;
            8'h2A : a[0:7] = 8'h54;
            8'h2B : a[0:7] = 8'h56;
            8'h2C : a[0:7] = 8'h58;
            8'h2D : a[0:7] = 8'h5A;
            8'h2E : a[0:7] = 8'h5C;
            8'h2F : a[0:7] = 8'h5E;
            8'h30 : a[0:7] = 8'h60;
            8'h31 : a[0:7] = 8'h62;
            8'h32 : a[0:7] = 8'h64;
            8'h33 : a[0:7] = 8'h66;
            8'h34 : a[0:7] = 8'h68;
            8'h35 : a[0:7] = 8'h6A;
            8'h36 : a[0:7] = 8'h6C;
            8'h37 : a[0:7] = 8'h6E;
            8'h38 : a[0:7] = 8'h70;
            8'h39 : a[0:7] = 8'h72;
            8'h3A : a[0:7] = 8'h74;
            8'h3B : a[0:7] = 8'h76;
            8'h3C : a[0:7] = 8'h78;
            8'h3D : a[0:7] = 8'h7A;
            8'h3E : a[0:7] = 8'h7C;
            8'h3F : a[0:7] = 8'h7E;
            8'h40 : a[0:7] = 8'h80;
            8'h41 : a[0:7] = 8'h82;
            8'h42 : a[0:7] = 8'h84;
            8'h43 : a[0:7] = 8'h86;
            8'h44 : a[0:7] = 8'h88;
            8'h45 : a[0:7] = 8'h8A;
            8'h46 : a[0:7] = 8'h8C;
            8'h47 : a[0:7] = 8'h8E;
            8'h48 : a[0:7] = 8'h90;
            8'h49 : a[0:7] = 8'h92;
            8'h4A : a[0:7] = 8'h94;
            8'h4B : a[0:7] = 8'h96;
            8'h4C : a[0:7] = 8'h98;
            8'h4D : a[0:7] = 8'h9A;
            8'h4E : a[0:7] = 8'h9C;
            8'h4F : a[0:7] = 8'h9E;
            8'h50 : a[0:7] = 8'hA0;
            8'h51 : a[0:7] = 8'hA2;
            8'h52 : a[0:7] = 8'hA4;
            8'h53 : a[0:7] = 8'hA6;
            8'h54 : a[0:7] = 8'hA8;
            8'h55 : a[0:7] = 8'hAA;
            8'h56 : a[0:7] = 8'hAC;
            8'h57 : a[0:7] = 8'hAE;
            8'h58 : a[0:7] = 8'hB0;
            8'h59 : a[0:7] = 8'hB2;
            8'h5A : a[0:7] = 8'hB4;
            8'h5B : a[0:7] = 8'hB6;
            8'h5C : a[0:7] = 8'hB8;
            8'h5D : a[0:7] = 8'hBA;
            8'h5E : a[0:7] = 8'hBC;
            8'h5F : a[0:7] = 8'hBE;
            8'h60 : a[0:7] = 8'hC0;
            8'h61 : a[0:7] = 8'hC2;
            8'h62 : a[0:7] = 8'hC4;
            8'h63 : a[0:7] = 8'hC6;
            8'h64 : a[0:7] = 8'hC8;
            8'h65 : a[0:7] = 8'hCA;
            8'h66 : a[0:7] = 8'hCC;
            8'h67 : a[0:7] = 8'hCE;
            8'h68 : a[0:7] = 8'hD0;
            8'h69 : a[0:7] = 8'hD2;
            8'h6A : a[0:7] = 8'hD4;
            8'h6B : a[0:7] = 8'hD6;
            8'h6C : a[0:7] = 8'hD8;
            8'h6D : a[0:7] = 8'hDA;
            8'h6E : a[0:7] = 8'hDC;
            8'h6F : a[0:7] = 8'hDE;
            8'h70 : a[0:7] = 8'hE0;
            8'h71 : a[0:7] = 8'hE2;
            8'h72 : a[0:7] = 8'hE4;
            8'h73 : a[0:7] = 8'hE6;
            8'h74 : a[0:7] = 8'hE8;
            8'h75 : a[0:7] = 8'hEA;
            8'h76 : a[0:7] = 8'hEC;
            8'h77 : a[0:7] = 8'hEE;
            8'h78 : a[0:7] = 8'hF0;
            8'h79 : a[0:7] = 8'hF2;
            8'h7A : a[0:7] = 8'hF4;
            8'h7B : a[0:7] = 8'hF6;
            8'h7C : a[0:7] = 8'hF8;
            8'h7D : a[0:7] = 8'hFA;
            8'h7E : a[0:7] = 8'hFC;
            8'h7F : a[0:7] = 8'hFE;
            8'h80 : a[0:7] = 8'h1B;
            8'h81 : a[0:7] = 8'h19;
            8'h82 : a[0:7] = 8'h1F;
            8'h83 : a[0:7] = 8'h1D;
            8'h84 : a[0:7] = 8'h13;
            8'h85 : a[0:7] = 8'h11;
            8'h86 : a[0:7] = 8'h17;
            8'h87 : a[0:7] = 8'h15;
            8'h88 : a[0:7] = 8'hB;
            8'h89 : a[0:7] = 8'h9;
            8'h8A : a[0:7] = 8'hF;
            8'h8B : a[0:7] = 8'hD;
            8'h8C : a[0:7] = 8'h3;
            8'h8D : a[0:7] = 8'h1;
            8'h8E : a[0:7] = 8'h7;
            8'h8F : a[0:7] = 8'h5;
            8'h90 : a[0:7] = 8'h3B;
            8'h91 : a[0:7] = 8'h39;
            8'h92 : a[0:7] = 8'h3F;
            8'h93 : a[0:7] = 8'h3D;
            8'h94 : a[0:7] = 8'h33;
            8'h95 : a[0:7] = 8'h31;
            8'h96 : a[0:7] = 8'h37;
            8'h97 : a[0:7] = 8'h35;
            8'h98 : a[0:7] = 8'h2B;
            8'h99 : a[0:7] = 8'h29;
            8'h9A : a[0:7] = 8'h2F;
            8'h9B : a[0:7] = 8'h2D;
            8'h9C : a[0:7] = 8'h23;
            8'h9D : a[0:7] = 8'h21;
            8'h9E : a[0:7] = 8'h27;
            8'h9F : a[0:7] = 8'h25;
            8'hA0 : a[0:7] = 8'h5B;
            8'hA1 : a[0:7] = 8'h59;
            8'hA2 : a[0:7] = 8'h5F;
            8'hA3 : a[0:7] = 8'h5D;
            8'hA4 : a[0:7] = 8'h53;
            8'hA5 : a[0:7] = 8'h51;
            8'hA6 : a[0:7] = 8'h57;
            8'hA7 : a[0:7] = 8'h55;
            8'hA8 : a[0:7] = 8'h4B;
            8'hA9 : a[0:7] = 8'h49;
            8'hAA : a[0:7] = 8'h4F;
            8'hAB : a[0:7] = 8'h4D;
            8'hAC : a[0:7] = 8'h43;
            8'hAD : a[0:7] = 8'h41;
            8'hAE : a[0:7] = 8'h47;
            8'hAF : a[0:7] = 8'h45;
            8'hB0 : a[0:7] = 8'h7B;
            8'hB1 : a[0:7] = 8'h79;
            8'hB2 : a[0:7] = 8'h7F;
            8'hB3 : a[0:7] = 8'h7D;
            8'hB4 : a[0:7] = 8'h73;
            8'hB5 : a[0:7] = 8'h71;
            8'hB6 : a[0:7] = 8'h77;
            8'hB7 : a[0:7] = 8'h75;
            8'hB8 : a[0:7] = 8'h6B;
            8'hB9 : a[0:7] = 8'h69;
            8'hBA : a[0:7] = 8'h6F;
            8'hBB : a[0:7] = 8'h6D;
            8'hBC : a[0:7] = 8'h63;
            8'hBD : a[0:7] = 8'h61;
            8'hBE : a[0:7] = 8'h67;
            8'hBF : a[0:7] = 8'h65;
            8'hC0 : a[0:7] = 8'h9B;
            8'hC1 : a[0:7] = 8'h99;
            8'hC2 : a[0:7] = 8'h9F;
            8'hC3 : a[0:7] = 8'h9D;
            8'hC4 : a[0:7] = 8'h93;
            8'hC5 : a[0:7] = 8'h91;
            8'hC6 : a[0:7] = 8'h97;
            8'hC7 : a[0:7] = 8'h95;
            8'hC8 : a[0:7] = 8'h8B;
            8'hC9 : a[0:7] = 8'h89;
            8'hCA : a[0:7] = 8'h8F;
            8'hCB : a[0:7] = 8'h8D;
            8'hCC : a[0:7] = 8'h83;
            8'hCD : a[0:7] = 8'h81;
            8'hCE : a[0:7] = 8'h87;
            8'hCF : a[0:7] = 8'h85;
            8'hD0 : a[0:7] = 8'hBB;
            8'hD1 : a[0:7] = 8'hB9;
            8'hD2 : a[0:7] = 8'hBF;
            8'hD3 : a[0:7] = 8'hBD;
            8'hD4 : a[0:7] = 8'hB3;
            8'hD5 : a[0:7] = 8'hB1;
            8'hD6 : a[0:7] = 8'hB7;
            8'hD7 : a[0:7] = 8'hB5;
            8'hD8 : a[0:7] = 8'hAB;
            8'hD9 : a[0:7] = 8'hA9;
            8'hDA : a[0:7] = 8'hAF;
            8'hDB : a[0:7] = 8'hAD;
            8'hDC : a[0:7] = 8'hA3;
            8'hDD : a[0:7] = 8'hA1;
            8'hDE : a[0:7] = 8'hA7;
            8'hDF : a[0:7] = 8'hA5;
            8'hE0 : a[0:7] = 8'hDB;
            8'hE1 : a[0:7] = 8'hD9;
            8'hE2 : a[0:7] = 8'hDF;
            8'hE3 : a[0:7] = 8'hDD;
            8'hE4 : a[0:7] = 8'hD3;
            8'hE5 : a[0:7] = 8'hD1;
            8'hE6 : a[0:7] = 8'hD7;
            8'hE7 : a[0:7] = 8'hD5;
            8'hE8 : a[0:7] = 8'hCB;
            8'hE9 : a[0:7] = 8'hC9;
            8'hEA : a[0:7] = 8'hCF;
            8'hEB : a[0:7] = 8'hCD;
            8'hEC : a[0:7] = 8'hC3;
            8'hED : a[0:7] = 8'hC1;
            8'hEE : a[0:7] = 8'hC7;
            8'hEF : a[0:7] = 8'hC5;
            8'hF0 : a[0:7] = 8'hFB;
            8'hF1 : a[0:7] = 8'hF9;
            8'hF2 : a[0:7] = 8'hFF;
            8'hF3 : a[0:7] = 8'hFD;
            8'hF4 : a[0:7] = 8'hF3;
            8'hF5 : a[0:7] = 8'hF1;
            8'hF6 : a[0:7] = 8'hF7;
            8'hF7 : a[0:7] = 8'hF5;
            8'hF8 : a[0:7] = 8'hEB;
            8'hF9 : a[0:7] = 8'hE9;
            8'hFA : a[0:7] = 8'hEF;
            8'hFB : a[0:7] = 8'hED;
            8'hFC : a[0:7] = 8'hE3;
            8'hFD : a[0:7] = 8'hE1;
            8'hFE : a[0:7] = 8'hE7;
            8'hFF : a[0:7] = 8'hE5;
        endcase
    end

    always @(row[24:31]) begin
        // Multiplication with 3
        case (row[24:31])
            8'h0 : b[0:7] = 8'h0;
            8'h1 : b[0:7] = 8'h3;
            8'h2 : b[0:7] = 8'h6;
            8'h3 : b[0:7] = 8'h5;
            8'h4 : b[0:7] = 8'hC;
            8'h5 : b[0:7] = 8'hF;
            8'h6 : b[0:7] = 8'hA;
            8'h7 : b[0:7] = 8'h9;
            8'h8 : b[0:7] = 8'h18;
            8'h9 : b[0:7] = 8'h1B;
            8'hA : b[0:7] = 8'h1E;
            8'hB : b[0:7] = 8'h1D;
            8'hC : b[0:7] = 8'h14;
            8'hD : b[0:7] = 8'h17;
            8'hE : b[0:7] = 8'h12;
            8'hF : b[0:7] = 8'h11;
            8'h10 : b[0:7] = 8'h30;
            8'h11 : b[0:7] = 8'h33;
            8'h12 : b[0:7] = 8'h36;
            8'h13 : b[0:7] = 8'h35;
            8'h14 : b[0:7] = 8'h3C;
            8'h15 : b[0:7] = 8'h3F;
            8'h16 : b[0:7] = 8'h3A;
            8'h17 : b[0:7] = 8'h39;
            8'h18 : b[0:7] = 8'h28;
            8'h19 : b[0:7] = 8'h2B;
            8'h1A : b[0:7] = 8'h2E;
            8'h1B : b[0:7] = 8'h2D;
            8'h1C : b[0:7] = 8'h24;
            8'h1D : b[0:7] = 8'h27;
            8'h1E : b[0:7] = 8'h22;
            8'h1F : b[0:7] = 8'h21;
            8'h20 : b[0:7] = 8'h60;
            8'h21 : b[0:7] = 8'h63;
            8'h22 : b[0:7] = 8'h66;
            8'h23 : b[0:7] = 8'h65;
            8'h24 : b[0:7] = 8'h6C;
            8'h25 : b[0:7] = 8'h6F;
            8'h26 : b[0:7] = 8'h6A;
            8'h27 : b[0:7] = 8'h69;
            8'h28 : b[0:7] = 8'h78;
            8'h29 : b[0:7] = 8'h7B;
            8'h2A : b[0:7] = 8'h7E;
            8'h2B : b[0:7] = 8'h7D;
            8'h2C : b[0:7] = 8'h74;
            8'h2D : b[0:7] = 8'h77;
            8'h2E : b[0:7] = 8'h72;
            8'h2F : b[0:7] = 8'h71;
            8'h30 : b[0:7] = 8'h50;
            8'h31 : b[0:7] = 8'h53;
            8'h32 : b[0:7] = 8'h56;
            8'h33 : b[0:7] = 8'h55;
            8'h34 : b[0:7] = 8'h5C;
            8'h35 : b[0:7] = 8'h5F;
            8'h36 : b[0:7] = 8'h5A;
            8'h37 : b[0:7] = 8'h59;
            8'h38 : b[0:7] = 8'h48;
            8'h39 : b[0:7] = 8'h4B;
            8'h3A : b[0:7] = 8'h4E;
            8'h3B : b[0:7] = 8'h4D;
            8'h3C : b[0:7] = 8'h44;
            8'h3D : b[0:7] = 8'h47;
            8'h3E : b[0:7] = 8'h42;
            8'h3F : b[0:7] = 8'h41;
            8'h40 : b[0:7] = 8'hC0;
            8'h41 : b[0:7] = 8'hC3;
            8'h42 : b[0:7] = 8'hC6;
            8'h43 : b[0:7] = 8'hC5;
            8'h44 : b[0:7] = 8'hCC;
            8'h45 : b[0:7] = 8'hCF;
            8'h46 : b[0:7] = 8'hCA;
            8'h47 : b[0:7] = 8'hC9;
            8'h48 : b[0:7] = 8'hD8;
            8'h49 : b[0:7] = 8'hDB;
            8'h4A : b[0:7] = 8'hDE;
            8'h4B : b[0:7] = 8'hDD;
            8'h4C : b[0:7] = 8'hD4;
            8'h4D : b[0:7] = 8'hD7;
            8'h4E : b[0:7] = 8'hD2;
            8'h4F : b[0:7] = 8'hD1;
            8'h50 : b[0:7] = 8'hF0;
            8'h51 : b[0:7] = 8'hF3;
            8'h52 : b[0:7] = 8'hF6;
            8'h53 : b[0:7] = 8'hF5;
            8'h54 : b[0:7] = 8'hFC;
            8'h55 : b[0:7] = 8'hFF;
            8'h56 : b[0:7] = 8'hFA;
            8'h57 : b[0:7] = 8'hF9;
            8'h58 : b[0:7] = 8'hE8;
            8'h59 : b[0:7] = 8'hEB;
            8'h5A : b[0:7] = 8'hEE;
            8'h5B : b[0:7] = 8'hED;
            8'h5C : b[0:7] = 8'hE4;
            8'h5D : b[0:7] = 8'hE7;
            8'h5E : b[0:7] = 8'hE2;
            8'h5F : b[0:7] = 8'hE1;
            8'h60 : b[0:7] = 8'hA0;
            8'h61 : b[0:7] = 8'hA3;
            8'h62 : b[0:7] = 8'hA6;
            8'h63 : b[0:7] = 8'hA5;
            8'h64 : b[0:7] = 8'hAC;
            8'h65 : b[0:7] = 8'hAF;
            8'h66 : b[0:7] = 8'hAA;
            8'h67 : b[0:7] = 8'hA9;
            8'h68 : b[0:7] = 8'hB8;
            8'h69 : b[0:7] = 8'hBB;
            8'h6A : b[0:7] = 8'hBE;
            8'h6B : b[0:7] = 8'hBD;
            8'h6C : b[0:7] = 8'hB4;
            8'h6D : b[0:7] = 8'hB7;
            8'h6E : b[0:7] = 8'hB2;
            8'h6F : b[0:7] = 8'hB1;
            8'h70 : b[0:7] = 8'h90;
            8'h71 : b[0:7] = 8'h93;
            8'h72 : b[0:7] = 8'h96;
            8'h73 : b[0:7] = 8'h95;
            8'h74 : b[0:7] = 8'h9C;
            8'h75 : b[0:7] = 8'h9F;
            8'h76 : b[0:7] = 8'h9A;
            8'h77 : b[0:7] = 8'h99;
            8'h78 : b[0:7] = 8'h88;
            8'h79 : b[0:7] = 8'h8B;
            8'h7A : b[0:7] = 8'h8E;
            8'h7B : b[0:7] = 8'h8D;
            8'h7C : b[0:7] = 8'h84;
            8'h7D : b[0:7] = 8'h87;
            8'h7E : b[0:7] = 8'h82;
            8'h7F : b[0:7] = 8'h81;
            8'h80 : b[0:7] = 8'h9B;
            8'h81 : b[0:7] = 8'h98;
            8'h82 : b[0:7] = 8'h9D;
            8'h83 : b[0:7] = 8'h9E;
            8'h84 : b[0:7] = 8'h97;
            8'h85 : b[0:7] = 8'h94;
            8'h86 : b[0:7] = 8'h91;
            8'h87 : b[0:7] = 8'h92;
            8'h88 : b[0:7] = 8'h83;
            8'h89 : b[0:7] = 8'h80;
            8'h8A : b[0:7] = 8'h85;
            8'h8B : b[0:7] = 8'h86;
            8'h8C : b[0:7] = 8'h8F;
            8'h8D : b[0:7] = 8'h8C;
            8'h8E : b[0:7] = 8'h89;
            8'h8F : b[0:7] = 8'h8A;
            8'h90 : b[0:7] = 8'hAB;
            8'h91 : b[0:7] = 8'hA8;
            8'h92 : b[0:7] = 8'hAD;
            8'h93 : b[0:7] = 8'hAE;
            8'h94 : b[0:7] = 8'hA7;
            8'h95 : b[0:7] = 8'hA4;
            8'h96 : b[0:7] = 8'hA1;
            8'h97 : b[0:7] = 8'hA2;
            8'h98 : b[0:7] = 8'hB3;
            8'h99 : b[0:7] = 8'hB0;
            8'h9A : b[0:7] = 8'hB5;
            8'h9B : b[0:7] = 8'hB6;
            8'h9C : b[0:7] = 8'hBF;
            8'h9D : b[0:7] = 8'hBC;
            8'h9E : b[0:7] = 8'hB9;
            8'h9F : b[0:7] = 8'hBA;
            8'hA0 : b[0:7] = 8'hFB;
            8'hA1 : b[0:7] = 8'hF8;
            8'hA2 : b[0:7] = 8'hFD;
            8'hA3 : b[0:7] = 8'hFE;
            8'hA4 : b[0:7] = 8'hF7;
            8'hA5 : b[0:7] = 8'hF4;
            8'hA6 : b[0:7] = 8'hF1;
            8'hA7 : b[0:7] = 8'hF2;
            8'hA8 : b[0:7] = 8'hE3;
            8'hA9 : b[0:7] = 8'hE0;
            8'hAA : b[0:7] = 8'hE5;
            8'hAB : b[0:7] = 8'hE6;
            8'hAC : b[0:7] = 8'hEF;
            8'hAD : b[0:7] = 8'hEC;
            8'hAE : b[0:7] = 8'hE9;
            8'hAF : b[0:7] = 8'hEA;
            8'hB0 : b[0:7] = 8'hCB;
            8'hB1 : b[0:7] = 8'hC8;
            8'hB2 : b[0:7] = 8'hCD;
            8'hB3 : b[0:7] = 8'hCE;
            8'hB4 : b[0:7] = 8'hC7;
            8'hB5 : b[0:7] = 8'hC4;
            8'hB6 : b[0:7] = 8'hC1;
            8'hB7 : b[0:7] = 8'hC2;
            8'hB8 : b[0:7] = 8'hD3;
            8'hB9 : b[0:7] = 8'hD0;
            8'hBA : b[0:7] = 8'hD5;
            8'hBB : b[0:7] = 8'hD6;
            8'hBC : b[0:7] = 8'hDF;
            8'hBD : b[0:7] = 8'hDC;
            8'hBE : b[0:7] = 8'hD9;
            8'hBF : b[0:7] = 8'hDA;
            8'hC0 : b[0:7] = 8'h5B;
            8'hC1 : b[0:7] = 8'h58;
            8'hC2 : b[0:7] = 8'h5D;
            8'hC3 : b[0:7] = 8'h5E;
            8'hC4 : b[0:7] = 8'h57;
            8'hC5 : b[0:7] = 8'h54;
            8'hC6 : b[0:7] = 8'h51;
            8'hC7 : b[0:7] = 8'h52;
            8'hC8 : b[0:7] = 8'h43;
            8'hC9 : b[0:7] = 8'h40;
            8'hCA : b[0:7] = 8'h45;
            8'hCB : b[0:7] = 8'h46;
            8'hCC : b[0:7] = 8'h4F;
            8'hCD : b[0:7] = 8'h4C;
            8'hCE : b[0:7] = 8'h49;
            8'hCF : b[0:7] = 8'h4A;
            8'hD0 : b[0:7] = 8'h6B;
            8'hD1 : b[0:7] = 8'h68;
            8'hD2 : b[0:7] = 8'h6D;
            8'hD3 : b[0:7] = 8'h6E;
            8'hD4 : b[0:7] = 8'h67;
            8'hD5 : b[0:7] = 8'h64;
            8'hD6 : b[0:7] = 8'h61;
            8'hD7 : b[0:7] = 8'h62;
            8'hD8 : b[0:7] = 8'h73;
            8'hD9 : b[0:7] = 8'h70;
            8'hDA : b[0:7] = 8'h75;
            8'hDB : b[0:7] = 8'h76;
            8'hDC : b[0:7] = 8'h7F;
            8'hDD : b[0:7] = 8'h7C;
            8'hDE : b[0:7] = 8'h79;
            8'hDF : b[0:7] = 8'h7A;
            8'hE0 : b[0:7] = 8'h3B;
            8'hE1 : b[0:7] = 8'h38;
            8'hE2 : b[0:7] = 8'h3D;
            8'hE3 : b[0:7] = 8'h3E;
            8'hE4 : b[0:7] = 8'h37;
            8'hE5 : b[0:7] = 8'h34;
            8'hE6 : b[0:7] = 8'h31;
            8'hE7 : b[0:7] = 8'h32;
            8'hE8 : b[0:7] = 8'h23;
            8'hE9 : b[0:7] = 8'h20;
            8'hEA : b[0:7] = 8'h25;
            8'hEB : b[0:7] = 8'h26;
            8'hEC : b[0:7] = 8'h2F;
            8'hED : b[0:7] = 8'h2C;
            8'hEE : b[0:7] = 8'h29;
            8'hEF : b[0:7] = 8'h2A;
            8'hF0 : b[0:7] = 8'hB;
            8'hF1 : b[0:7] = 8'h8;
            8'hF2 : b[0:7] = 8'hD;
            8'hF3 : b[0:7] = 8'hE;
            8'hF4 : b[0:7] = 8'h7;
            8'hF5 : b[0:7] = 8'h4;
            8'hF6 : b[0:7] = 8'h1;
            8'hF7 : b[0:7] = 8'h2;
            8'hF8 : b[0:7] = 8'h13;
            8'hF9 : b[0:7] = 8'h10;
            8'hFA : b[0:7] = 8'h15;
            8'hFB : b[0:7] = 8'h16;
            8'hFC : b[0:7] = 8'h1F;
            8'hFD : b[0:7] = 8'h1C;
            8'hFE : b[0:7] = 8'h19;
            8'hFF : b[0:7] = 8'h1A;
        endcase
    end

    // Multiplication with 1
    always @(row[0:7]) begin
        c[0:7] = row[0:7];
    end

    // Multiplication with 1
    always @( row[8:15]) begin
        d[0:7] =  row[8:15];
    end

    assign output_row = a ^ b ^ c ^ d;
    
endmodule


module MixColumn4Row (
    input wire [0:31] row,
    output wire [0:7] output_row
);
    reg [0:7] a, b, c, d;

    // Multiplication with 2
    always @(row[24:31]) begin
        case (row[24:31])
            8'h0 : a[0:7] = 8'h0;
            8'h1 : a[0:7] = 8'h2;
            8'h2 : a[0:7] = 8'h4;
            8'h3 : a[0:7] = 8'h6;
            8'h4 : a[0:7] = 8'h8;
            8'h5 : a[0:7] = 8'hA;
            8'h6 : a[0:7] = 8'hC;
            8'h7 : a[0:7] = 8'hE;
            8'h8 : a[0:7] = 8'h10;
            8'h9 : a[0:7] = 8'h12;
            8'hA : a[0:7] = 8'h14;
            8'hB : a[0:7] = 8'h16;
            8'hC : a[0:7] = 8'h18;
            8'hD : a[0:7] = 8'h1A;
            8'hE : a[0:7] = 8'h1C;
            8'hF : a[0:7] = 8'h1E;
            8'h10 : a[0:7] = 8'h20;
            8'h11 : a[0:7] = 8'h22;
            8'h12 : a[0:7] = 8'h24;
            8'h13 : a[0:7] = 8'h26;
            8'h14 : a[0:7] = 8'h28;
            8'h15 : a[0:7] = 8'h2A;
            8'h16 : a[0:7] = 8'h2C;
            8'h17 : a[0:7] = 8'h2E;
            8'h18 : a[0:7] = 8'h30;
            8'h19 : a[0:7] = 8'h32;
            8'h1A : a[0:7] = 8'h34;
            8'h1B : a[0:7] = 8'h36;
            8'h1C : a[0:7] = 8'h38;
            8'h1D : a[0:7] = 8'h3A;
            8'h1E : a[0:7] = 8'h3C;
            8'h1F : a[0:7] = 8'h3E;
            8'h20 : a[0:7] = 8'h40;
            8'h21 : a[0:7] = 8'h42;
            8'h22 : a[0:7] = 8'h44;
            8'h23 : a[0:7] = 8'h46;
            8'h24 : a[0:7] = 8'h48;
            8'h25 : a[0:7] = 8'h4A;
            8'h26 : a[0:7] = 8'h4C;
            8'h27 : a[0:7] = 8'h4E;
            8'h28 : a[0:7] = 8'h50;
            8'h29 : a[0:7] = 8'h52;
            8'h2A : a[0:7] = 8'h54;
            8'h2B : a[0:7] = 8'h56;
            8'h2C : a[0:7] = 8'h58;
            8'h2D : a[0:7] = 8'h5A;
            8'h2E : a[0:7] = 8'h5C;
            8'h2F : a[0:7] = 8'h5E;
            8'h30 : a[0:7] = 8'h60;
            8'h31 : a[0:7] = 8'h62;
            8'h32 : a[0:7] = 8'h64;
            8'h33 : a[0:7] = 8'h66;
            8'h34 : a[0:7] = 8'h68;
            8'h35 : a[0:7] = 8'h6A;
            8'h36 : a[0:7] = 8'h6C;
            8'h37 : a[0:7] = 8'h6E;
            8'h38 : a[0:7] = 8'h70;
            8'h39 : a[0:7] = 8'h72;
            8'h3A : a[0:7] = 8'h74;
            8'h3B : a[0:7] = 8'h76;
            8'h3C : a[0:7] = 8'h78;
            8'h3D : a[0:7] = 8'h7A;
            8'h3E : a[0:7] = 8'h7C;
            8'h3F : a[0:7] = 8'h7E;
            8'h40 : a[0:7] = 8'h80;
            8'h41 : a[0:7] = 8'h82;
            8'h42 : a[0:7] = 8'h84;
            8'h43 : a[0:7] = 8'h86;
            8'h44 : a[0:7] = 8'h88;
            8'h45 : a[0:7] = 8'h8A;
            8'h46 : a[0:7] = 8'h8C;
            8'h47 : a[0:7] = 8'h8E;
            8'h48 : a[0:7] = 8'h90;
            8'h49 : a[0:7] = 8'h92;
            8'h4A : a[0:7] = 8'h94;
            8'h4B : a[0:7] = 8'h96;
            8'h4C : a[0:7] = 8'h98;
            8'h4D : a[0:7] = 8'h9A;
            8'h4E : a[0:7] = 8'h9C;
            8'h4F : a[0:7] = 8'h9E;
            8'h50 : a[0:7] = 8'hA0;
            8'h51 : a[0:7] = 8'hA2;
            8'h52 : a[0:7] = 8'hA4;
            8'h53 : a[0:7] = 8'hA6;
            8'h54 : a[0:7] = 8'hA8;
            8'h55 : a[0:7] = 8'hAA;
            8'h56 : a[0:7] = 8'hAC;
            8'h57 : a[0:7] = 8'hAE;
            8'h58 : a[0:7] = 8'hB0;
            8'h59 : a[0:7] = 8'hB2;
            8'h5A : a[0:7] = 8'hB4;
            8'h5B : a[0:7] = 8'hB6;
            8'h5C : a[0:7] = 8'hB8;
            8'h5D : a[0:7] = 8'hBA;
            8'h5E : a[0:7] = 8'hBC;
            8'h5F : a[0:7] = 8'hBE;
            8'h60 : a[0:7] = 8'hC0;
            8'h61 : a[0:7] = 8'hC2;
            8'h62 : a[0:7] = 8'hC4;
            8'h63 : a[0:7] = 8'hC6;
            8'h64 : a[0:7] = 8'hC8;
            8'h65 : a[0:7] = 8'hCA;
            8'h66 : a[0:7] = 8'hCC;
            8'h67 : a[0:7] = 8'hCE;
            8'h68 : a[0:7] = 8'hD0;
            8'h69 : a[0:7] = 8'hD2;
            8'h6A : a[0:7] = 8'hD4;
            8'h6B : a[0:7] = 8'hD6;
            8'h6C : a[0:7] = 8'hD8;
            8'h6D : a[0:7] = 8'hDA;
            8'h6E : a[0:7] = 8'hDC;
            8'h6F : a[0:7] = 8'hDE;
            8'h70 : a[0:7] = 8'hE0;
            8'h71 : a[0:7] = 8'hE2;
            8'h72 : a[0:7] = 8'hE4;
            8'h73 : a[0:7] = 8'hE6;
            8'h74 : a[0:7] = 8'hE8;
            8'h75 : a[0:7] = 8'hEA;
            8'h76 : a[0:7] = 8'hEC;
            8'h77 : a[0:7] = 8'hEE;
            8'h78 : a[0:7] = 8'hF0;
            8'h79 : a[0:7] = 8'hF2;
            8'h7A : a[0:7] = 8'hF4;
            8'h7B : a[0:7] = 8'hF6;
            8'h7C : a[0:7] = 8'hF8;
            8'h7D : a[0:7] = 8'hFA;
            8'h7E : a[0:7] = 8'hFC;
            8'h7F : a[0:7] = 8'hFE;
            8'h80 : a[0:7] = 8'h1B;
            8'h81 : a[0:7] = 8'h19;
            8'h82 : a[0:7] = 8'h1F;
            8'h83 : a[0:7] = 8'h1D;
            8'h84 : a[0:7] = 8'h13;
            8'h85 : a[0:7] = 8'h11;
            8'h86 : a[0:7] = 8'h17;
            8'h87 : a[0:7] = 8'h15;
            8'h88 : a[0:7] = 8'hB;
            8'h89 : a[0:7] = 8'h9;
            8'h8A : a[0:7] = 8'hF;
            8'h8B : a[0:7] = 8'hD;
            8'h8C : a[0:7] = 8'h3;
            8'h8D : a[0:7] = 8'h1;
            8'h8E : a[0:7] = 8'h7;
            8'h8F : a[0:7] = 8'h5;
            8'h90 : a[0:7] = 8'h3B;
            8'h91 : a[0:7] = 8'h39;
            8'h92 : a[0:7] = 8'h3F;
            8'h93 : a[0:7] = 8'h3D;
            8'h94 : a[0:7] = 8'h33;
            8'h95 : a[0:7] = 8'h31;
            8'h96 : a[0:7] = 8'h37;
            8'h97 : a[0:7] = 8'h35;
            8'h98 : a[0:7] = 8'h2B;
            8'h99 : a[0:7] = 8'h29;
            8'h9A : a[0:7] = 8'h2F;
            8'h9B : a[0:7] = 8'h2D;
            8'h9C : a[0:7] = 8'h23;
            8'h9D : a[0:7] = 8'h21;
            8'h9E : a[0:7] = 8'h27;
            8'h9F : a[0:7] = 8'h25;
            8'hA0 : a[0:7] = 8'h5B;
            8'hA1 : a[0:7] = 8'h59;
            8'hA2 : a[0:7] = 8'h5F;
            8'hA3 : a[0:7] = 8'h5D;
            8'hA4 : a[0:7] = 8'h53;
            8'hA5 : a[0:7] = 8'h51;
            8'hA6 : a[0:7] = 8'h57;
            8'hA7 : a[0:7] = 8'h55;
            8'hA8 : a[0:7] = 8'h4B;
            8'hA9 : a[0:7] = 8'h49;
            8'hAA : a[0:7] = 8'h4F;
            8'hAB : a[0:7] = 8'h4D;
            8'hAC : a[0:7] = 8'h43;
            8'hAD : a[0:7] = 8'h41;
            8'hAE : a[0:7] = 8'h47;
            8'hAF : a[0:7] = 8'h45;
            8'hB0 : a[0:7] = 8'h7B;
            8'hB1 : a[0:7] = 8'h79;
            8'hB2 : a[0:7] = 8'h7F;
            8'hB3 : a[0:7] = 8'h7D;
            8'hB4 : a[0:7] = 8'h73;
            8'hB5 : a[0:7] = 8'h71;
            8'hB6 : a[0:7] = 8'h77;
            8'hB7 : a[0:7] = 8'h75;
            8'hB8 : a[0:7] = 8'h6B;
            8'hB9 : a[0:7] = 8'h69;
            8'hBA : a[0:7] = 8'h6F;
            8'hBB : a[0:7] = 8'h6D;
            8'hBC : a[0:7] = 8'h63;
            8'hBD : a[0:7] = 8'h61;
            8'hBE : a[0:7] = 8'h67;
            8'hBF : a[0:7] = 8'h65;
            8'hC0 : a[0:7] = 8'h9B;
            8'hC1 : a[0:7] = 8'h99;
            8'hC2 : a[0:7] = 8'h9F;
            8'hC3 : a[0:7] = 8'h9D;
            8'hC4 : a[0:7] = 8'h93;
            8'hC5 : a[0:7] = 8'h91;
            8'hC6 : a[0:7] = 8'h97;
            8'hC7 : a[0:7] = 8'h95;
            8'hC8 : a[0:7] = 8'h8B;
            8'hC9 : a[0:7] = 8'h89;
            8'hCA : a[0:7] = 8'h8F;
            8'hCB : a[0:7] = 8'h8D;
            8'hCC : a[0:7] = 8'h83;
            8'hCD : a[0:7] = 8'h81;
            8'hCE : a[0:7] = 8'h87;
            8'hCF : a[0:7] = 8'h85;
            8'hD0 : a[0:7] = 8'hBB;
            8'hD1 : a[0:7] = 8'hB9;
            8'hD2 : a[0:7] = 8'hBF;
            8'hD3 : a[0:7] = 8'hBD;
            8'hD4 : a[0:7] = 8'hB3;
            8'hD5 : a[0:7] = 8'hB1;
            8'hD6 : a[0:7] = 8'hB7;
            8'hD7 : a[0:7] = 8'hB5;
            8'hD8 : a[0:7] = 8'hAB;
            8'hD9 : a[0:7] = 8'hA9;
            8'hDA : a[0:7] = 8'hAF;
            8'hDB : a[0:7] = 8'hAD;
            8'hDC : a[0:7] = 8'hA3;
            8'hDD : a[0:7] = 8'hA1;
            8'hDE : a[0:7] = 8'hA7;
            8'hDF : a[0:7] = 8'hA5;
            8'hE0 : a[0:7] = 8'hDB;
            8'hE1 : a[0:7] = 8'hD9;
            8'hE2 : a[0:7] = 8'hDF;
            8'hE3 : a[0:7] = 8'hDD;
            8'hE4 : a[0:7] = 8'hD3;
            8'hE5 : a[0:7] = 8'hD1;
            8'hE6 : a[0:7] = 8'hD7;
            8'hE7 : a[0:7] = 8'hD5;
            8'hE8 : a[0:7] = 8'hCB;
            8'hE9 : a[0:7] = 8'hC9;
            8'hEA : a[0:7] = 8'hCF;
            8'hEB : a[0:7] = 8'hCD;
            8'hEC : a[0:7] = 8'hC3;
            8'hED : a[0:7] = 8'hC1;
            8'hEE : a[0:7] = 8'hC7;
            8'hEF : a[0:7] = 8'hC5;
            8'hF0 : a[0:7] = 8'hFB;
            8'hF1 : a[0:7] = 8'hF9;
            8'hF2 : a[0:7] = 8'hFF;
            8'hF3 : a[0:7] = 8'hFD;
            8'hF4 : a[0:7] = 8'hF3;
            8'hF5 : a[0:7] = 8'hF1;
            8'hF6 : a[0:7] = 8'hF7;
            8'hF7 : a[0:7] = 8'hF5;
            8'hF8 : a[0:7] = 8'hEB;
            8'hF9 : a[0:7] = 8'hE9;
            8'hFA : a[0:7] = 8'hEF;
            8'hFB : a[0:7] = 8'hED;
            8'hFC : a[0:7] = 8'hE3;
            8'hFD : a[0:7] = 8'hE1;
            8'hFE : a[0:7] = 8'hE7;
            8'hFF : a[0:7] = 8'hE5;
        endcase
    end

    always @(row[0:7]) begin
        // Multiplication with 3
        case (row[0:7])
            8'h0 : b[0:7] = 8'h0;
            8'h1 : b[0:7] = 8'h3;
            8'h2 : b[0:7] = 8'h6;
            8'h3 : b[0:7] = 8'h5;
            8'h4 : b[0:7] = 8'hC;
            8'h5 : b[0:7] = 8'hF;
            8'h6 : b[0:7] = 8'hA;
            8'h7 : b[0:7] = 8'h9;
            8'h8 : b[0:7] = 8'h18;
            8'h9 : b[0:7] = 8'h1B;
            8'hA : b[0:7] = 8'h1E;
            8'hB : b[0:7] = 8'h1D;
            8'hC : b[0:7] = 8'h14;
            8'hD : b[0:7] = 8'h17;
            8'hE : b[0:7] = 8'h12;
            8'hF : b[0:7] = 8'h11;
            8'h10 : b[0:7] = 8'h30;
            8'h11 : b[0:7] = 8'h33;
            8'h12 : b[0:7] = 8'h36;
            8'h13 : b[0:7] = 8'h35;
            8'h14 : b[0:7] = 8'h3C;
            8'h15 : b[0:7] = 8'h3F;
            8'h16 : b[0:7] = 8'h3A;
            8'h17 : b[0:7] = 8'h39;
            8'h18 : b[0:7] = 8'h28;
            8'h19 : b[0:7] = 8'h2B;
            8'h1A : b[0:7] = 8'h2E;
            8'h1B : b[0:7] = 8'h2D;
            8'h1C : b[0:7] = 8'h24;
            8'h1D : b[0:7] = 8'h27;
            8'h1E : b[0:7] = 8'h22;
            8'h1F : b[0:7] = 8'h21;
            8'h20 : b[0:7] = 8'h60;
            8'h21 : b[0:7] = 8'h63;
            8'h22 : b[0:7] = 8'h66;
            8'h23 : b[0:7] = 8'h65;
            8'h24 : b[0:7] = 8'h6C;
            8'h25 : b[0:7] = 8'h6F;
            8'h26 : b[0:7] = 8'h6A;
            8'h27 : b[0:7] = 8'h69;
            8'h28 : b[0:7] = 8'h78;
            8'h29 : b[0:7] = 8'h7B;
            8'h2A : b[0:7] = 8'h7E;
            8'h2B : b[0:7] = 8'h7D;
            8'h2C : b[0:7] = 8'h74;
            8'h2D : b[0:7] = 8'h77;
            8'h2E : b[0:7] = 8'h72;
            8'h2F : b[0:7] = 8'h71;
            8'h30 : b[0:7] = 8'h50;
            8'h31 : b[0:7] = 8'h53;
            8'h32 : b[0:7] = 8'h56;
            8'h33 : b[0:7] = 8'h55;
            8'h34 : b[0:7] = 8'h5C;
            8'h35 : b[0:7] = 8'h5F;
            8'h36 : b[0:7] = 8'h5A;
            8'h37 : b[0:7] = 8'h59;
            8'h38 : b[0:7] = 8'h48;
            8'h39 : b[0:7] = 8'h4B;
            8'h3A : b[0:7] = 8'h4E;
            8'h3B : b[0:7] = 8'h4D;
            8'h3C : b[0:7] = 8'h44;
            8'h3D : b[0:7] = 8'h47;
            8'h3E : b[0:7] = 8'h42;
            8'h3F : b[0:7] = 8'h41;
            8'h40 : b[0:7] = 8'hC0;
            8'h41 : b[0:7] = 8'hC3;
            8'h42 : b[0:7] = 8'hC6;
            8'h43 : b[0:7] = 8'hC5;
            8'h44 : b[0:7] = 8'hCC;
            8'h45 : b[0:7] = 8'hCF;
            8'h46 : b[0:7] = 8'hCA;
            8'h47 : b[0:7] = 8'hC9;
            8'h48 : b[0:7] = 8'hD8;
            8'h49 : b[0:7] = 8'hDB;
            8'h4A : b[0:7] = 8'hDE;
            8'h4B : b[0:7] = 8'hDD;
            8'h4C : b[0:7] = 8'hD4;
            8'h4D : b[0:7] = 8'hD7;
            8'h4E : b[0:7] = 8'hD2;
            8'h4F : b[0:7] = 8'hD1;
            8'h50 : b[0:7] = 8'hF0;
            8'h51 : b[0:7] = 8'hF3;
            8'h52 : b[0:7] = 8'hF6;
            8'h53 : b[0:7] = 8'hF5;
            8'h54 : b[0:7] = 8'hFC;
            8'h55 : b[0:7] = 8'hFF;
            8'h56 : b[0:7] = 8'hFA;
            8'h57 : b[0:7] = 8'hF9;
            8'h58 : b[0:7] = 8'hE8;
            8'h59 : b[0:7] = 8'hEB;
            8'h5A : b[0:7] = 8'hEE;
            8'h5B : b[0:7] = 8'hED;
            8'h5C : b[0:7] = 8'hE4;
            8'h5D : b[0:7] = 8'hE7;
            8'h5E : b[0:7] = 8'hE2;
            8'h5F : b[0:7] = 8'hE1;
            8'h60 : b[0:7] = 8'hA0;
            8'h61 : b[0:7] = 8'hA3;
            8'h62 : b[0:7] = 8'hA6;
            8'h63 : b[0:7] = 8'hA5;
            8'h64 : b[0:7] = 8'hAC;
            8'h65 : b[0:7] = 8'hAF;
            8'h66 : b[0:7] = 8'hAA;
            8'h67 : b[0:7] = 8'hA9;
            8'h68 : b[0:7] = 8'hB8;
            8'h69 : b[0:7] = 8'hBB;
            8'h6A : b[0:7] = 8'hBE;
            8'h6B : b[0:7] = 8'hBD;
            8'h6C : b[0:7] = 8'hB4;
            8'h6D : b[0:7] = 8'hB7;
            8'h6E : b[0:7] = 8'hB2;
            8'h6F : b[0:7] = 8'hB1;
            8'h70 : b[0:7] = 8'h90;
            8'h71 : b[0:7] = 8'h93;
            8'h72 : b[0:7] = 8'h96;
            8'h73 : b[0:7] = 8'h95;
            8'h74 : b[0:7] = 8'h9C;
            8'h75 : b[0:7] = 8'h9F;
            8'h76 : b[0:7] = 8'h9A;
            8'h77 : b[0:7] = 8'h99;
            8'h78 : b[0:7] = 8'h88;
            8'h79 : b[0:7] = 8'h8B;
            8'h7A : b[0:7] = 8'h8E;
            8'h7B : b[0:7] = 8'h8D;
            8'h7C : b[0:7] = 8'h84;
            8'h7D : b[0:7] = 8'h87;
            8'h7E : b[0:7] = 8'h82;
            8'h7F : b[0:7] = 8'h81;
            8'h80 : b[0:7] = 8'h9B;
            8'h81 : b[0:7] = 8'h98;
            8'h82 : b[0:7] = 8'h9D;
            8'h83 : b[0:7] = 8'h9E;
            8'h84 : b[0:7] = 8'h97;
            8'h85 : b[0:7] = 8'h94;
            8'h86 : b[0:7] = 8'h91;
            8'h87 : b[0:7] = 8'h92;
            8'h88 : b[0:7] = 8'h83;
            8'h89 : b[0:7] = 8'h80;
            8'h8A : b[0:7] = 8'h85;
            8'h8B : b[0:7] = 8'h86;
            8'h8C : b[0:7] = 8'h8F;
            8'h8D : b[0:7] = 8'h8C;
            8'h8E : b[0:7] = 8'h89;
            8'h8F : b[0:7] = 8'h8A;
            8'h90 : b[0:7] = 8'hAB;
            8'h91 : b[0:7] = 8'hA8;
            8'h92 : b[0:7] = 8'hAD;
            8'h93 : b[0:7] = 8'hAE;
            8'h94 : b[0:7] = 8'hA7;
            8'h95 : b[0:7] = 8'hA4;
            8'h96 : b[0:7] = 8'hA1;
            8'h97 : b[0:7] = 8'hA2;
            8'h98 : b[0:7] = 8'hB3;
            8'h99 : b[0:7] = 8'hB0;
            8'h9A : b[0:7] = 8'hB5;
            8'h9B : b[0:7] = 8'hB6;
            8'h9C : b[0:7] = 8'hBF;
            8'h9D : b[0:7] = 8'hBC;
            8'h9E : b[0:7] = 8'hB9;
            8'h9F : b[0:7] = 8'hBA;
            8'hA0 : b[0:7] = 8'hFB;
            8'hA1 : b[0:7] = 8'hF8;
            8'hA2 : b[0:7] = 8'hFD;
            8'hA3 : b[0:7] = 8'hFE;
            8'hA4 : b[0:7] = 8'hF7;
            8'hA5 : b[0:7] = 8'hF4;
            8'hA6 : b[0:7] = 8'hF1;
            8'hA7 : b[0:7] = 8'hF2;
            8'hA8 : b[0:7] = 8'hE3;
            8'hA9 : b[0:7] = 8'hE0;
            8'hAA : b[0:7] = 8'hE5;
            8'hAB : b[0:7] = 8'hE6;
            8'hAC : b[0:7] = 8'hEF;
            8'hAD : b[0:7] = 8'hEC;
            8'hAE : b[0:7] = 8'hE9;
            8'hAF : b[0:7] = 8'hEA;
            8'hB0 : b[0:7] = 8'hCB;
            8'hB1 : b[0:7] = 8'hC8;
            8'hB2 : b[0:7] = 8'hCD;
            8'hB3 : b[0:7] = 8'hCE;
            8'hB4 : b[0:7] = 8'hC7;
            8'hB5 : b[0:7] = 8'hC4;
            8'hB6 : b[0:7] = 8'hC1;
            8'hB7 : b[0:7] = 8'hC2;
            8'hB8 : b[0:7] = 8'hD3;
            8'hB9 : b[0:7] = 8'hD0;
            8'hBA : b[0:7] = 8'hD5;
            8'hBB : b[0:7] = 8'hD6;
            8'hBC : b[0:7] = 8'hDF;
            8'hBD : b[0:7] = 8'hDC;
            8'hBE : b[0:7] = 8'hD9;
            8'hBF : b[0:7] = 8'hDA;
            8'hC0 : b[0:7] = 8'h5B;
            8'hC1 : b[0:7] = 8'h58;
            8'hC2 : b[0:7] = 8'h5D;
            8'hC3 : b[0:7] = 8'h5E;
            8'hC4 : b[0:7] = 8'h57;
            8'hC5 : b[0:7] = 8'h54;
            8'hC6 : b[0:7] = 8'h51;
            8'hC7 : b[0:7] = 8'h52;
            8'hC8 : b[0:7] = 8'h43;
            8'hC9 : b[0:7] = 8'h40;
            8'hCA : b[0:7] = 8'h45;
            8'hCB : b[0:7] = 8'h46;
            8'hCC : b[0:7] = 8'h4F;
            8'hCD : b[0:7] = 8'h4C;
            8'hCE : b[0:7] = 8'h49;
            8'hCF : b[0:7] = 8'h4A;
            8'hD0 : b[0:7] = 8'h6B;
            8'hD1 : b[0:7] = 8'h68;
            8'hD2 : b[0:7] = 8'h6D;
            8'hD3 : b[0:7] = 8'h6E;
            8'hD4 : b[0:7] = 8'h67;
            8'hD5 : b[0:7] = 8'h64;
            8'hD6 : b[0:7] = 8'h61;
            8'hD7 : b[0:7] = 8'h62;
            8'hD8 : b[0:7] = 8'h73;
            8'hD9 : b[0:7] = 8'h70;
            8'hDA : b[0:7] = 8'h75;
            8'hDB : b[0:7] = 8'h76;
            8'hDC : b[0:7] = 8'h7F;
            8'hDD : b[0:7] = 8'h7C;
            8'hDE : b[0:7] = 8'h79;
            8'hDF : b[0:7] = 8'h7A;
            8'hE0 : b[0:7] = 8'h3B;
            8'hE1 : b[0:7] = 8'h38;
            8'hE2 : b[0:7] = 8'h3D;
            8'hE3 : b[0:7] = 8'h3E;
            8'hE4 : b[0:7] = 8'h37;
            8'hE5 : b[0:7] = 8'h34;
            8'hE6 : b[0:7] = 8'h31;
            8'hE7 : b[0:7] = 8'h32;
            8'hE8 : b[0:7] = 8'h23;
            8'hE9 : b[0:7] = 8'h20;
            8'hEA : b[0:7] = 8'h25;
            8'hEB : b[0:7] = 8'h26;
            8'hEC : b[0:7] = 8'h2F;
            8'hED : b[0:7] = 8'h2C;
            8'hEE : b[0:7] = 8'h29;
            8'hEF : b[0:7] = 8'h2A;
            8'hF0 : b[0:7] = 8'hB;
            8'hF1 : b[0:7] = 8'h8;
            8'hF2 : b[0:7] = 8'hD;
            8'hF3 : b[0:7] = 8'hE;
            8'hF4 : b[0:7] = 8'h7;
            8'hF5 : b[0:7] = 8'h4;
            8'hF6 : b[0:7] = 8'h1;
            8'hF7 : b[0:7] = 8'h2;
            8'hF8 : b[0:7] = 8'h13;
            8'hF9 : b[0:7] = 8'h10;
            8'hFA : b[0:7] = 8'h15;
            8'hFB : b[0:7] = 8'h16;
            8'hFC : b[0:7] = 8'h1F;
            8'hFD : b[0:7] = 8'h1C;
            8'hFE : b[0:7] = 8'h19;
            8'hFF : b[0:7] = 8'h1A;
        endcase
    end

    // Multiplication with 1
    always @(row[8:15]) begin
        c[0:7] = row[8:15];
    end

    // Multiplication with 1
    always @(row[16:23]) begin
        d[0:7] = row[16:23];
    end

    assign output_row = a ^ b ^ c ^ d;
    
endmodule


module MixColumn (
    input wire [0:31] row,
    output wire [0:31] output_row
);
    wire [0:7] a, b, c, d;

    MixColumn1Row MixColumn1RowModule(row[0:31], a[0:7]);
    MixColumn2Row MixColumn2RowModule(row[0:31], b[0:7]);
    MixColumn3Row MixColumn3RowModule(row[0:31], c[0:7]);
    MixColumn4Row MixColumn4RowModule(row[0:31], d[0:7]);

    assign output_row[0:7] = a[0:7];
    assign output_row[8:15] = b[0:7];
    assign output_row[16:23] = c[0:7];
    assign output_row[24:31] = d[0:7];
    

    
endmodule